-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_0_start: Boolean;
  signal convTranspose_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_ConvTranspose_input_pipe_734_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_734_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_734_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_716_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_734_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_1 : boolean;
  signal addr_of_475_final_reg_ack_1 : boolean;
  signal type_cast_689_inst_req_0 : boolean;
  signal addr_of_475_final_reg_req_1 : boolean;
  signal type_cast_513_inst_ack_1 : boolean;
  signal type_cast_513_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_478_inst_req_0 : boolean;
  signal type_cast_513_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_478_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_478_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_478_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 : boolean;
  signal type_cast_513_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1044_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_685_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_685_inst_req_0 : boolean;
  signal if_stmt_625_branch_ack_0 : boolean;
  signal type_cast_31_inst_req_0 : boolean;
  signal type_cast_31_inst_ack_0 : boolean;
  signal type_cast_31_inst_req_1 : boolean;
  signal type_cast_567_inst_ack_0 : boolean;
  signal type_cast_31_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_509_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_1 : boolean;
  signal type_cast_567_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 : boolean;
  signal type_cast_531_inst_ack_1 : boolean;
  signal type_cast_44_inst_req_0 : boolean;
  signal type_cast_44_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1044_inst_ack_0 : boolean;
  signal type_cast_44_inst_req_1 : boolean;
  signal type_cast_44_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_52_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_52_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_509_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_52_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_52_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_509_inst_req_0 : boolean;
  signal type_cast_531_inst_req_1 : boolean;
  signal if_stmt_625_branch_ack_1 : boolean;
  signal type_cast_56_inst_req_0 : boolean;
  signal type_cast_56_inst_ack_0 : boolean;
  signal type_cast_56_inst_req_1 : boolean;
  signal type_cast_56_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_152_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_152_inst_ack_1 : boolean;
  signal if_stmt_1369_branch_ack_1 : boolean;
  signal type_cast_585_inst_req_0 : boolean;
  signal type_cast_1247_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_998_inst_req_1 : boolean;
  signal type_cast_1049_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1004_inst_req_0 : boolean;
  signal type_cast_69_inst_req_0 : boolean;
  signal type_cast_69_inst_ack_0 : boolean;
  signal type_cast_69_inst_req_1 : boolean;
  signal type_cast_69_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_ack_0 : boolean;
  signal type_cast_1042_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_77_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_77_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_509_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_77_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_77_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1004_inst_ack_0 : boolean;
  signal type_cast_81_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1007_inst_req_0 : boolean;
  signal type_cast_81_inst_ack_0 : boolean;
  signal type_cast_81_inst_req_1 : boolean;
  signal type_cast_81_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1054_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1004_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_0 : boolean;
  signal type_cast_531_inst_ack_0 : boolean;
  signal type_cast_94_inst_req_0 : boolean;
  signal type_cast_94_inst_ack_0 : boolean;
  signal type_cast_94_inst_req_1 : boolean;
  signal type_cast_94_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1044_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_102_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_102_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_102_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_102_inst_ack_1 : boolean;
  signal type_cast_702_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_0 : boolean;
  signal addr_of_682_final_reg_ack_1 : boolean;
  signal type_cast_531_inst_req_0 : boolean;
  signal type_cast_106_inst_req_0 : boolean;
  signal type_cast_106_inst_ack_0 : boolean;
  signal type_cast_106_inst_req_1 : boolean;
  signal type_cast_106_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 : boolean;
  signal type_cast_702_inst_req_1 : boolean;
  signal addr_of_682_final_reg_req_1 : boolean;
  signal if_stmt_625_branch_req_0 : boolean;
  signal WPIPE_Block0_start_998_inst_ack_1 : boolean;
  signal type_cast_585_inst_ack_1 : boolean;
  signal type_cast_119_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_1 : boolean;
  signal type_cast_119_inst_ack_0 : boolean;
  signal type_cast_119_inst_req_1 : boolean;
  signal type_cast_119_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_127_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_127_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_127_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_563_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_127_inst_ack_1 : boolean;
  signal addr_of_682_final_reg_ack_0 : boolean;
  signal WPIPE_Block2_start_1072_inst_req_1 : boolean;
  signal type_cast_585_inst_req_1 : boolean;
  signal type_cast_131_inst_req_0 : boolean;
  signal type_cast_131_inst_ack_0 : boolean;
  signal type_cast_131_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_563_inst_req_1 : boolean;
  signal type_cast_131_inst_ack_1 : boolean;
  signal type_cast_720_inst_ack_1 : boolean;
  signal type_cast_495_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 : boolean;
  signal type_cast_495_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 : boolean;
  signal addr_of_682_final_reg_req_0 : boolean;
  signal type_cast_603_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_998_inst_req_0 : boolean;
  signal type_cast_144_inst_req_0 : boolean;
  signal type_cast_144_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_1 : boolean;
  signal type_cast_144_inst_req_1 : boolean;
  signal type_cast_144_inst_ack_1 : boolean;
  signal type_cast_720_inst_req_1 : boolean;
  signal type_cast_585_inst_ack_0 : boolean;
  signal type_cast_603_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1044_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_152_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_563_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_152_inst_ack_0 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_545_inst_ack_1 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal type_cast_482_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_545_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 : boolean;
  signal type_cast_482_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 : boolean;
  signal type_cast_156_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_563_inst_req_0 : boolean;
  signal type_cast_156_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_998_inst_ack_0 : boolean;
  signal type_cast_156_inst_req_1 : boolean;
  signal type_cast_156_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_0 : boolean;
  signal type_cast_1312_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 : boolean;
  signal type_cast_495_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 : boolean;
  signal type_cast_702_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_1 : boolean;
  signal type_cast_1049_inst_ack_1 : boolean;
  signal type_cast_169_inst_req_0 : boolean;
  signal type_cast_169_inst_ack_0 : boolean;
  signal ptr_deref_611_store_0_ack_1 : boolean;
  signal type_cast_169_inst_req_1 : boolean;
  signal type_cast_169_inst_ack_1 : boolean;
  signal type_cast_495_inst_req_0 : boolean;
  signal type_cast_603_inst_ack_0 : boolean;
  signal type_cast_603_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_177_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_177_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_177_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_177_inst_ack_1 : boolean;
  signal type_cast_181_inst_req_0 : boolean;
  signal type_cast_181_inst_ack_0 : boolean;
  signal ptr_deref_611_store_0_req_1 : boolean;
  signal type_cast_181_inst_req_1 : boolean;
  signal type_cast_181_inst_ack_1 : boolean;
  signal type_cast_720_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 : boolean;
  signal type_cast_702_inst_req_0 : boolean;
  signal type_cast_194_inst_req_0 : boolean;
  signal type_cast_194_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_1 : boolean;
  signal type_cast_194_inst_ack_1 : boolean;
  signal type_cast_720_inst_req_0 : boolean;
  signal type_cast_203_inst_req_0 : boolean;
  signal type_cast_203_inst_ack_0 : boolean;
  signal type_cast_203_inst_req_1 : boolean;
  signal type_cast_203_inst_ack_1 : boolean;
  signal type_cast_652_inst_ack_1 : boolean;
  signal type_cast_207_inst_req_0 : boolean;
  signal type_cast_207_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_0 : boolean;
  signal type_cast_207_inst_req_1 : boolean;
  signal type_cast_207_inst_ack_1 : boolean;
  signal type_cast_652_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_0 : boolean;
  signal ptr_deref_611_store_0_ack_0 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal ptr_deref_611_store_0_req_0 : boolean;
  signal type_cast_248_inst_req_0 : boolean;
  signal type_cast_549_inst_ack_1 : boolean;
  signal type_cast_248_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_0 : boolean;
  signal type_cast_248_inst_req_1 : boolean;
  signal type_cast_549_inst_req_1 : boolean;
  signal type_cast_248_inst_ack_1 : boolean;
  signal type_cast_652_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_req_1 : boolean;
  signal type_cast_252_inst_req_0 : boolean;
  signal type_cast_252_inst_ack_0 : boolean;
  signal type_cast_252_inst_req_1 : boolean;
  signal type_cast_252_inst_ack_1 : boolean;
  signal type_cast_652_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_req_0 : boolean;
  signal type_cast_256_inst_req_0 : boolean;
  signal type_cast_256_inst_ack_0 : boolean;
  signal type_cast_256_inst_req_1 : boolean;
  signal type_cast_549_inst_ack_0 : boolean;
  signal type_cast_256_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1054_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_ack_0 : boolean;
  signal type_cast_260_inst_req_0 : boolean;
  signal type_cast_549_inst_req_0 : boolean;
  signal type_cast_260_inst_ack_0 : boolean;
  signal type_cast_260_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1069_inst_req_1 : boolean;
  signal type_cast_260_inst_ack_1 : boolean;
  signal phi_stmt_669_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_1 : boolean;
  signal type_cast_282_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1343_inst_ack_0 : boolean;
  signal type_cast_282_inst_ack_0 : boolean;
  signal type_cast_282_inst_req_1 : boolean;
  signal type_cast_282_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 : boolean;
  signal array_obj_ref_681_index_offset_ack_1 : boolean;
  signal type_cast_295_inst_req_0 : boolean;
  signal type_cast_295_inst_ack_0 : boolean;
  signal type_cast_295_inst_req_1 : boolean;
  signal type_cast_295_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_ack_1 : boolean;
  signal array_obj_ref_681_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_1 : boolean;
  signal type_cast_307_inst_req_0 : boolean;
  signal type_cast_307_inst_ack_0 : boolean;
  signal type_cast_307_inst_req_1 : boolean;
  signal type_cast_307_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 : boolean;
  signal array_obj_ref_681_index_offset_ack_0 : boolean;
  signal type_cast_320_inst_req_0 : boolean;
  signal type_cast_320_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_1 : boolean;
  signal type_cast_320_inst_ack_1 : boolean;
  signal type_cast_689_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_716_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_ack_1 : boolean;
  signal array_obj_ref_681_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_685_inst_ack_1 : boolean;
  signal type_cast_332_inst_req_0 : boolean;
  signal type_cast_332_inst_ack_0 : boolean;
  signal type_cast_332_inst_req_1 : boolean;
  signal type_cast_332_inst_ack_1 : boolean;
  signal type_cast_689_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_716_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_1 : boolean;
  signal type_cast_1049_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_685_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1004_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_527_inst_ack_1 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_1049_inst_ack_0 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_ack_1 : boolean;
  signal type_cast_1042_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_527_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_1 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_716_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_378_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_378_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_378_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1007_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_378_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_527_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_527_inst_req_0 : boolean;
  signal type_cast_382_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_545_inst_ack_0 : boolean;
  signal type_cast_382_inst_ack_0 : boolean;
  signal type_cast_382_inst_req_1 : boolean;
  signal type_cast_382_inst_ack_1 : boolean;
  signal type_cast_689_inst_ack_0 : boolean;
  signal type_cast_482_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_545_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 : boolean;
  signal type_cast_482_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 : boolean;
  signal type_cast_567_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_1 : boolean;
  signal type_cast_395_inst_req_0 : boolean;
  signal type_cast_395_inst_ack_0 : boolean;
  signal type_cast_395_inst_req_1 : boolean;
  signal type_cast_395_inst_ack_1 : boolean;
  signal type_cast_1105_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal if_stmt_409_branch_req_0 : boolean;
  signal if_stmt_409_branch_ack_1 : boolean;
  signal if_stmt_409_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_1 : boolean;
  signal type_cast_567_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_1 : boolean;
  signal if_stmt_424_branch_req_0 : boolean;
  signal if_stmt_424_branch_ack_1 : boolean;
  signal if_stmt_424_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_1 : boolean;
  signal type_cast_445_inst_req_0 : boolean;
  signal type_cast_445_inst_ack_0 : boolean;
  signal type_cast_445_inst_req_1 : boolean;
  signal type_cast_445_inst_ack_1 : boolean;
  signal array_obj_ref_474_index_offset_req_0 : boolean;
  signal array_obj_ref_474_index_offset_ack_0 : boolean;
  signal array_obj_ref_474_index_offset_req_1 : boolean;
  signal array_obj_ref_474_index_offset_ack_1 : boolean;
  signal addr_of_475_final_reg_req_0 : boolean;
  signal addr_of_475_final_reg_ack_0 : boolean;
  signal type_cast_738_inst_req_0 : boolean;
  signal type_cast_738_inst_ack_0 : boolean;
  signal type_cast_738_inst_req_1 : boolean;
  signal type_cast_738_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_0 : boolean;
  signal if_stmt_1369_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_752_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_752_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1010_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_752_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1066_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_752_inst_ack_1 : boolean;
  signal type_cast_1098_inst_ack_1 : boolean;
  signal type_cast_1098_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_ack_0 : boolean;
  signal type_cast_1042_inst_ack_0 : boolean;
  signal type_cast_756_inst_req_0 : boolean;
  signal type_cast_756_inst_ack_0 : boolean;
  signal type_cast_756_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1066_inst_req_1 : boolean;
  signal type_cast_756_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1100_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1010_inst_req_1 : boolean;
  signal phi_stmt_913_req_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_770_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_770_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_770_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_770_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_req_0 : boolean;
  signal type_cast_1042_inst_req_0 : boolean;
  signal phi_stmt_669_req_1 : boolean;
  signal type_cast_774_inst_req_0 : boolean;
  signal type_cast_774_inst_ack_0 : boolean;
  signal type_cast_774_inst_req_1 : boolean;
  signal type_cast_774_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1100_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1066_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1010_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_ack_1 : boolean;
  signal type_cast_1098_inst_ack_0 : boolean;
  signal type_cast_1098_inst_req_0 : boolean;
  signal type_cast_1312_inst_ack_0 : boolean;
  signal type_cast_792_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1066_inst_req_0 : boolean;
  signal type_cast_792_inst_ack_0 : boolean;
  signal type_cast_792_inst_req_1 : boolean;
  signal type_cast_792_inst_ack_1 : boolean;
  signal type_cast_1312_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_806_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_806_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1010_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_806_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_806_inst_ack_1 : boolean;
  signal if_stmt_1369_branch_ack_0 : boolean;
  signal type_cast_810_inst_req_0 : boolean;
  signal type_cast_810_inst_ack_0 : boolean;
  signal type_cast_810_inst_req_1 : boolean;
  signal type_cast_810_inst_ack_1 : boolean;
  signal phi_stmt_1241_ack_0 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1063_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal ptr_deref_818_store_0_req_0 : boolean;
  signal ptr_deref_818_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal ptr_deref_818_store_0_req_1 : boolean;
  signal ptr_deref_818_store_0_ack_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_0 : boolean;
  signal type_cast_1312_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1054_inst_ack_0 : boolean;
  signal if_stmt_832_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1054_inst_req_0 : boolean;
  signal if_stmt_832_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_1001_inst_ack_1 : boolean;
  signal if_stmt_832_branch_ack_0 : boolean;
  signal type_cast_843_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1063_inst_req_1 : boolean;
  signal type_cast_843_inst_ack_0 : boolean;
  signal type_cast_843_inst_req_1 : boolean;
  signal type_cast_843_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1100_inst_ack_0 : boolean;
  signal type_cast_1105_inst_ack_1 : boolean;
  signal type_cast_847_inst_req_0 : boolean;
  signal type_cast_847_inst_ack_0 : boolean;
  signal type_cast_847_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1063_inst_ack_0 : boolean;
  signal type_cast_847_inst_ack_1 : boolean;
  signal type_cast_1105_inst_req_1 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1063_inst_req_0 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_1 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1100_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1001_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_1 : boolean;
  signal if_stmt_869_branch_req_0 : boolean;
  signal if_stmt_869_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_1001_inst_ack_0 : boolean;
  signal if_stmt_869_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1051_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1051_inst_req_1 : boolean;
  signal type_cast_916_inst_req_0 : boolean;
  signal type_cast_896_inst_req_0 : boolean;
  signal type_cast_896_inst_ack_0 : boolean;
  signal type_cast_896_inst_req_1 : boolean;
  signal type_cast_896_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1001_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_0 : boolean;
  signal array_obj_ref_925_index_offset_req_0 : boolean;
  signal array_obj_ref_925_index_offset_ack_0 : boolean;
  signal array_obj_ref_925_index_offset_req_1 : boolean;
  signal array_obj_ref_925_index_offset_ack_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1343_inst_req_0 : boolean;
  signal addr_of_926_final_reg_req_0 : boolean;
  signal addr_of_926_final_reg_ack_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_0 : boolean;
  signal addr_of_926_final_reg_req_1 : boolean;
  signal addr_of_926_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1069_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1060_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1007_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_0 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal ptr_deref_929_store_0_req_0 : boolean;
  signal ptr_deref_929_store_0_ack_0 : boolean;
  signal WPIPE_Block0_start_994_inst_req_1 : boolean;
  signal ptr_deref_929_store_0_req_1 : boolean;
  signal ptr_deref_929_store_0_ack_1 : boolean;
  signal WPIPE_Block1_start_1007_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_0 : boolean;
  signal if_stmt_944_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal if_stmt_944_branch_ack_1 : boolean;
  signal if_stmt_944_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1051_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1051_inst_req_0 : boolean;
  signal type_cast_1105_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_954_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_954_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_954_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_954_inst_ack_1 : boolean;
  signal type_cast_1332_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_958_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_958_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1343_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_958_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_958_inst_ack_1 : boolean;
  signal phi_stmt_1241_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1343_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_963_inst_req_0 : boolean;
  signal WPIPE_Block0_start_963_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_963_inst_req_1 : boolean;
  signal WPIPE_Block0_start_963_inst_ack_1 : boolean;
  signal type_cast_1332_inst_ack_0 : boolean;
  signal type_cast_1322_inst_req_0 : boolean;
  signal WPIPE_Block0_start_966_inst_req_0 : boolean;
  signal WPIPE_Block0_start_966_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_966_inst_req_1 : boolean;
  signal WPIPE_Block0_start_966_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_969_inst_req_0 : boolean;
  signal WPIPE_Block0_start_969_inst_ack_0 : boolean;
  signal type_cast_916_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_969_inst_req_1 : boolean;
  signal WPIPE_Block0_start_969_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_972_inst_req_0 : boolean;
  signal WPIPE_Block0_start_972_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_972_inst_req_1 : boolean;
  signal WPIPE_Block0_start_972_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_975_inst_req_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_req_1 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_1 : boolean;
  signal type_cast_1322_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_978_inst_req_0 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_978_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_req_0 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_981_inst_req_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_984_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_1 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_987_inst_req_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_req_1 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_req_0 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_req_0 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1340_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1107_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1107_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1107_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1107_inst_ack_1 : boolean;
  signal type_cast_1322_inst_ack_1 : boolean;
  signal type_cast_1322_inst_req_1 : boolean;
  signal type_cast_1247_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1110_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1110_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1340_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1110_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1110_inst_ack_1 : boolean;
  signal phi_stmt_669_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_1 : boolean;
  signal type_cast_1247_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_req_1 : boolean;
  signal type_cast_672_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_1 : boolean;
  signal type_cast_1247_inst_req_0 : boolean;
  signal type_cast_672_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1119_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1119_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1340_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1119_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1119_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1122_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1122_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1340_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1122_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1122_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_req_1 : boolean;
  signal phi_stmt_462_ack_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1128_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1128_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1128_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1128_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_0 : boolean;
  signal phi_stmt_462_req_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_1 : boolean;
  signal type_cast_468_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1337_inst_ack_1 : boolean;
  signal phi_stmt_1241_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_0 : boolean;
  signal type_cast_468_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1337_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_1 : boolean;
  signal type_cast_468_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1337_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_0 : boolean;
  signal type_cast_468_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1337_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_1 : boolean;
  signal type_cast_1154_inst_req_0 : boolean;
  signal type_cast_1154_inst_ack_0 : boolean;
  signal type_cast_1154_inst_req_1 : boolean;
  signal type_cast_1154_inst_ack_1 : boolean;
  signal type_cast_672_inst_ack_0 : boolean;
  signal type_cast_672_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1156_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1156_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1156_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1156_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1334_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1349_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1349_inst_req_1 : boolean;
  signal type_cast_1161_inst_req_0 : boolean;
  signal type_cast_1161_inst_ack_0 : boolean;
  signal type_cast_1161_inst_req_1 : boolean;
  signal type_cast_1161_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1334_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1349_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1349_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1163_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1163_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1163_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1163_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1334_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1166_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1166_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1166_inst_req_1 : boolean;
  signal phi_stmt_462_req_0 : boolean;
  signal WPIPE_Block3_start_1166_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1334_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1346_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1346_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1176_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1176_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1176_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1176_inst_ack_1 : boolean;
  signal phi_stmt_913_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1346_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1179_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1179_inst_ack_0 : boolean;
  signal type_cast_1332_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1179_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1179_inst_ack_1 : boolean;
  signal type_cast_1332_inst_req_1 : boolean;
  signal phi_stmt_913_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1346_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1182_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1182_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1182_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1182_inst_ack_1 : boolean;
  signal type_cast_916_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1185_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1185_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1185_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1185_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_ack_1 : boolean;
  signal if_stmt_1197_branch_req_0 : boolean;
  signal if_stmt_1197_branch_ack_1 : boolean;
  signal if_stmt_1197_branch_ack_0 : boolean;
  signal type_cast_1224_inst_req_0 : boolean;
  signal type_cast_1224_inst_ack_0 : boolean;
  signal type_cast_1224_inst_req_1 : boolean;
  signal type_cast_1224_inst_ack_1 : boolean;
  signal array_obj_ref_1253_index_offset_req_0 : boolean;
  signal array_obj_ref_1253_index_offset_ack_0 : boolean;
  signal array_obj_ref_1253_index_offset_req_1 : boolean;
  signal array_obj_ref_1253_index_offset_ack_1 : boolean;
  signal addr_of_1254_final_reg_req_0 : boolean;
  signal addr_of_1254_final_reg_ack_0 : boolean;
  signal addr_of_1254_final_reg_req_1 : boolean;
  signal addr_of_1254_final_reg_ack_1 : boolean;
  signal ptr_deref_1258_load_0_req_0 : boolean;
  signal ptr_deref_1258_load_0_ack_0 : boolean;
  signal ptr_deref_1258_load_0_req_1 : boolean;
  signal ptr_deref_1258_load_0_ack_1 : boolean;
  signal type_cast_1262_inst_req_0 : boolean;
  signal type_cast_1262_inst_ack_0 : boolean;
  signal type_cast_1262_inst_req_1 : boolean;
  signal type_cast_1262_inst_ack_1 : boolean;
  signal type_cast_1272_inst_req_0 : boolean;
  signal type_cast_1272_inst_ack_0 : boolean;
  signal type_cast_1272_inst_req_1 : boolean;
  signal type_cast_1272_inst_ack_1 : boolean;
  signal type_cast_1282_inst_req_0 : boolean;
  signal type_cast_1282_inst_ack_0 : boolean;
  signal type_cast_1282_inst_req_1 : boolean;
  signal type_cast_1282_inst_ack_1 : boolean;
  signal type_cast_1292_inst_req_0 : boolean;
  signal type_cast_1292_inst_ack_0 : boolean;
  signal type_cast_1292_inst_req_1 : boolean;
  signal type_cast_1292_inst_ack_1 : boolean;
  signal type_cast_1302_inst_req_0 : boolean;
  signal type_cast_1302_inst_ack_0 : boolean;
  signal type_cast_1302_inst_req_1 : boolean;
  signal type_cast_1302_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_0: Block -- control-path 
    signal convTranspose_CP_0_elements: BooleanArray(457 downto 0);
    -- 
  begin -- 
    convTranspose_CP_0_elements(0) <= convTranspose_CP_0_start;
    convTranspose_CP_0_symbol <= convTranspose_CP_0_elements(457);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_25/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/branch_block_stmt_25__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Update/cr
      -- 
    rr_96_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_96_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_27_inst_req_0); -- 
    cr_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_31_inst_req_1); -- 
    cr_143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_44_inst_req_1); -- 
    cr_171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_56_inst_req_1); -- 
    cr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_69_inst_req_1); -- 
    cr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_81_inst_req_1); -- 
    cr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_94_inst_req_1); -- 
    cr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_106_inst_req_1); -- 
    cr_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_119_inst_req_1); -- 
    cr_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_131_inst_req_1); -- 
    cr_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_144_inst_req_1); -- 
    cr_773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_357_inst_req_1); -- 
    cr_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_156_inst_req_1); -- 
    cr_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_169_inst_req_1); -- 
    cr_451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_181_inst_req_1); -- 
    cr_479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_194_inst_req_1); -- 
    cr_493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_203_inst_req_1); -- 
    cr_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_207_inst_req_1); -- 
    cr_521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_211_inst_req_1); -- 
    cr_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_248_inst_req_1); -- 
    cr_549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_252_inst_req_1); -- 
    cr_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_256_inst_req_1); -- 
    cr_577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_260_inst_req_1); -- 
    cr_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_282_inst_req_1); -- 
    cr_633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_295_inst_req_1); -- 
    cr_661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_307_inst_req_1); -- 
    cr_689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_320_inst_req_1); -- 
    cr_717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_332_inst_req_1); -- 
    cr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_345_inst_req_1); -- 
    cr_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_370_inst_req_1); -- 
    cr_829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_382_inst_req_1); -- 
    cr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(0), ack => type_cast_395_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_update_start_
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Update/cr
      -- 
    ra_97_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_27_inst_ack_0, ack => convTranspose_CP_0_elements(1)); -- 
    cr_101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_27_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_27_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Sample/rr
      -- 
    ca_102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_27_inst_ack_1, ack => convTranspose_CP_0_elements(2)); -- 
    rr_110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(2), ack => type_cast_31_inst_req_0); -- 
    rr_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Sample/ra
      -- 
    ra_111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_31_inst_ack_0, ack => convTranspose_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_31_Update/ca
      -- 
    ca_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_31_inst_ack_1, ack => convTranspose_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_update_start_
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Update/cr
      -- 
    ra_125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_0, ack => convTranspose_CP_0_elements(5)); -- 
    cr_129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(5), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_40_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Sample/rr
      -- 
    ca_130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_1, ack => convTranspose_CP_0_elements(6)); -- 
    rr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(6), ack => type_cast_44_inst_req_0); -- 
    rr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(6), ack => RPIPE_ConvTranspose_input_pipe_52_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Sample/ra
      -- 
    ra_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_0, ack => convTranspose_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_44_Update/ca
      -- 
    ca_144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_1, ack => convTranspose_CP_0_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_update_start_
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Update/cr
      -- 
    ra_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_52_inst_ack_0, ack => convTranspose_CP_0_elements(9)); -- 
    cr_157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(9), ack => RPIPE_ConvTranspose_input_pipe_52_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_52_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_sample_start_
      -- 
    ca_158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_52_inst_ack_1, ack => convTranspose_CP_0_elements(10)); -- 
    rr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(10), ack => type_cast_56_inst_req_0); -- 
    rr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(10), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Sample/ra
      -- 
    ra_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_56_inst_ack_0, ack => convTranspose_CP_0_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_56_Update/ca
      -- 
    ca_172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_56_inst_ack_1, ack => convTranspose_CP_0_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_update_start_
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Update/cr
      -- 
    ra_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_0, ack => convTranspose_CP_0_elements(13)); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(13), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_65_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_1, ack => convTranspose_CP_0_elements(14)); -- 
    rr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(14), ack => type_cast_69_inst_req_0); -- 
    rr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(14), ack => RPIPE_ConvTranspose_input_pipe_77_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Sample/ra
      -- 
    ra_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_0, ack => convTranspose_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_69_Update/ca
      -- 
    ca_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_1, ack => convTranspose_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_update_start_
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Update/cr
      -- 
    ra_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_77_inst_ack_0, ack => convTranspose_CP_0_elements(17)); -- 
    cr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(17), ack => RPIPE_ConvTranspose_input_pipe_77_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_77_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Sample/rr
      -- 
    ca_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_77_inst_ack_1, ack => convTranspose_CP_0_elements(18)); -- 
    rr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(18), ack => type_cast_81_inst_req_0); -- 
    rr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(18), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Sample/ra
      -- 
    ra_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_81_inst_ack_0, ack => convTranspose_CP_0_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_81_Update/ca
      -- 
    ca_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_81_inst_ack_1, ack => convTranspose_CP_0_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_update_start_
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Update/cr
      -- 
    ra_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_0, ack => convTranspose_CP_0_elements(21)); -- 
    cr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(21), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_90_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Sample/rr
      -- 
    ca_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_1, ack => convTranspose_CP_0_elements(22)); -- 
    rr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(22), ack => type_cast_94_inst_req_0); -- 
    rr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(22), ack => RPIPE_ConvTranspose_input_pipe_102_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Sample/ra
      -- 
    ra_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_0, ack => convTranspose_CP_0_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_94_Update/ca
      -- 
    ca_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_1, ack => convTranspose_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_update_start_
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Update/cr
      -- 
    ra_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_102_inst_ack_0, ack => convTranspose_CP_0_elements(25)); -- 
    cr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(25), ack => RPIPE_ConvTranspose_input_pipe_102_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_102_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Sample/rr
      -- 
    ca_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_102_inst_ack_1, ack => convTranspose_CP_0_elements(26)); -- 
    rr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(26), ack => type_cast_106_inst_req_0); -- 
    rr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(26), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Sample/ra
      -- 
    ra_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_106_inst_ack_0, ack => convTranspose_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_106_Update/ca
      -- 
    ca_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_106_inst_ack_1, ack => convTranspose_CP_0_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_update_start_
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Update/cr
      -- 
    ra_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_0, ack => convTranspose_CP_0_elements(29)); -- 
    cr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(29), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_115_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Sample/rr
      -- 
    ca_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_1, ack => convTranspose_CP_0_elements(30)); -- 
    rr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(30), ack => type_cast_119_inst_req_0); -- 
    rr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(30), ack => RPIPE_ConvTranspose_input_pipe_127_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Sample/ra
      -- 
    ra_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_0, ack => convTranspose_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_119_Update/ca
      -- 
    ca_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_1, ack => convTranspose_CP_0_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_update_start_
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Update/cr
      -- 
    ra_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_127_inst_ack_0, ack => convTranspose_CP_0_elements(33)); -- 
    cr_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(33), ack => RPIPE_ConvTranspose_input_pipe_127_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_127_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Sample/rr
      -- 
    ca_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_127_inst_ack_1, ack => convTranspose_CP_0_elements(34)); -- 
    rr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(34), ack => type_cast_131_inst_req_0); -- 
    rr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(34), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Sample/ra
      -- 
    ra_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_131_inst_ack_0, ack => convTranspose_CP_0_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_131_Update/ca
      -- 
    ca_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_131_inst_ack_1, ack => convTranspose_CP_0_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_update_start_
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Update/cr
      -- 
    ra_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_0, ack => convTranspose_CP_0_elements(37)); -- 
    cr_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(37), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_140_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Sample/rr
      -- 
    ca_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_1, ack => convTranspose_CP_0_elements(38)); -- 
    rr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(38), ack => RPIPE_ConvTranspose_input_pipe_152_inst_req_0); -- 
    rr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(38), ack => type_cast_144_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Sample/ra
      -- 
    ra_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_0, ack => convTranspose_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_144_Update/ca
      -- 
    ca_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_1, ack => convTranspose_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_update_start_
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Sample/ra
      -- 
    ra_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_152_inst_ack_0, ack => convTranspose_CP_0_elements(41)); -- 
    cr_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(41), ack => RPIPE_ConvTranspose_input_pipe_152_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_152_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Sample/rr
      -- 
    ca_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_152_inst_ack_1, ack => convTranspose_CP_0_elements(42)); -- 
    rr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(42), ack => type_cast_156_inst_req_0); -- 
    rr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(42), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Sample/ra
      -- 
    ra_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_156_inst_ack_0, ack => convTranspose_CP_0_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_156_Update/ca
      -- 
    ca_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_156_inst_ack_1, ack => convTranspose_CP_0_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_update_start_
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Update/cr
      -- 
    ra_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_0, ack => convTranspose_CP_0_elements(45)); -- 
    cr_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(45), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_165_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Sample/rr
      -- 
    ca_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_1, ack => convTranspose_CP_0_elements(46)); -- 
    rr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(46), ack => RPIPE_ConvTranspose_input_pipe_177_inst_req_0); -- 
    rr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(46), ack => type_cast_169_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Sample/ra
      -- 
    ra_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_0, ack => convTranspose_CP_0_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_169_Update/ca
      -- 
    ca_424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_1, ack => convTranspose_CP_0_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_update_start_
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Update/cr
      -- 
    ra_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_177_inst_ack_0, ack => convTranspose_CP_0_elements(49)); -- 
    cr_437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(49), ack => RPIPE_ConvTranspose_input_pipe_177_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_177_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Sample/rr
      -- 
    ca_438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_177_inst_ack_1, ack => convTranspose_CP_0_elements(50)); -- 
    rr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(50), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_0); -- 
    rr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(50), ack => type_cast_181_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Sample/ra
      -- 
    ra_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_0, ack => convTranspose_CP_0_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_181_Update/ca
      -- 
    ca_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_1, ack => convTranspose_CP_0_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_update_start_
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Update/cr
      -- 
    ra_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_0, ack => convTranspose_CP_0_elements(53)); -- 
    cr_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(53), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	78 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_190_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Sample/rr
      -- 
    ca_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_1, ack => convTranspose_CP_0_elements(54)); -- 
    rr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(54), ack => RPIPE_ConvTranspose_input_pipe_278_inst_req_0); -- 
    rr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(54), ack => type_cast_194_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Sample/ra
      -- 
    ra_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_0, ack => convTranspose_CP_0_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_194_Update/ca
      -- 
    ca_480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_1, ack => convTranspose_CP_0_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Sample/rr
      -- 
    rr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(57), ack => type_cast_203_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(4) & convTranspose_CP_0_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Sample/ra
      -- 
    ra_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_203_inst_ack_0, ack => convTranspose_CP_0_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_203_Update/ca
      -- 
    ca_494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_203_inst_ack_1, ack => convTranspose_CP_0_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Sample/rr
      -- 
    rr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(60), ack => type_cast_207_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(12) & convTranspose_CP_0_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Sample/ra
      -- 
    ra_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_0, ack => convTranspose_CP_0_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_207_Update/ca
      -- 
    ca_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_1, ack => convTranspose_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Sample/rr
      -- 
    rr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(63), ack => type_cast_211_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(20) & convTranspose_CP_0_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Sample/ra
      -- 
    ra_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => convTranspose_CP_0_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_211_Update/ca
      -- 
    ca_522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => convTranspose_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Sample/rr
      -- 
    rr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(66), ack => type_cast_248_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(28) & convTranspose_CP_0_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Sample/ra
      -- 
    ra_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_248_inst_ack_0, ack => convTranspose_CP_0_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_248_Update/ca
      -- 
    ca_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_248_inst_ack_1, ack => convTranspose_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Sample/rr
      -- 
    rr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(69), ack => type_cast_252_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(40) & convTranspose_CP_0_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Sample/ra
      -- 
    ra_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_252_inst_ack_0, ack => convTranspose_CP_0_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_252_Update/ca
      -- 
    ca_550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_252_inst_ack_1, ack => convTranspose_CP_0_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Sample/rr
      -- 
    rr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(72), ack => type_cast_256_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(44) & convTranspose_CP_0_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Sample/ra
      -- 
    ra_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_0, ack => convTranspose_CP_0_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_256_Update/ca
      -- 
    ca_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_1, ack => convTranspose_CP_0_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Sample/rr
      -- 
    rr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(75), ack => type_cast_260_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(52) & convTranspose_CP_0_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Sample/ra
      -- 
    ra_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_0, ack => convTranspose_CP_0_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_260_Update/ca
      -- 
    ca_578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_1, ack => convTranspose_CP_0_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_update_start_
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Update/cr
      -- 
    ra_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_278_inst_ack_0, ack => convTranspose_CP_0_elements(78)); -- 
    cr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(78), ack => RPIPE_ConvTranspose_input_pipe_278_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_278_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Sample/rr
      -- 
    ca_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_278_inst_ack_1, ack => convTranspose_CP_0_elements(79)); -- 
    rr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(79), ack => type_cast_282_inst_req_0); -- 
    rr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(79), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Sample/ra
      -- 
    ra_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_0, ack => convTranspose_CP_0_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_282_Update/ca
      -- 
    ca_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_1, ack => convTranspose_CP_0_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_update_start_
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Update/cr
      -- 
    ra_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_0, ack => convTranspose_CP_0_elements(82)); -- 
    cr_619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(82), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_291_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Sample/rr
      -- 
    ca_620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_1, ack => convTranspose_CP_0_elements(83)); -- 
    rr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(83), ack => type_cast_295_inst_req_0); -- 
    rr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(83), ack => RPIPE_ConvTranspose_input_pipe_303_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Sample/ra
      -- 
    ra_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_0, ack => convTranspose_CP_0_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_295_Update/ca
      -- 
    ca_634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_1, ack => convTranspose_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_update_start_
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Update/cr
      -- 
    ra_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_303_inst_ack_0, ack => convTranspose_CP_0_elements(86)); -- 
    cr_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(86), ack => RPIPE_ConvTranspose_input_pipe_303_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_303_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Sample/rr
      -- 
    ca_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_303_inst_ack_1, ack => convTranspose_CP_0_elements(87)); -- 
    rr_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(87), ack => type_cast_307_inst_req_0); -- 
    rr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(87), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Sample/ra
      -- 
    ra_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_307_inst_ack_0, ack => convTranspose_CP_0_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_307_Update/ca
      -- 
    ca_662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_307_inst_ack_1, ack => convTranspose_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_update_start_
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Update/cr
      -- 
    ra_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_0, ack => convTranspose_CP_0_elements(90)); -- 
    cr_675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(90), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_316_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Sample/rr
      -- 
    ca_676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_1, ack => convTranspose_CP_0_elements(91)); -- 
    rr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(91), ack => type_cast_320_inst_req_0); -- 
    rr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(91), ack => RPIPE_ConvTranspose_input_pipe_328_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Sample/ra
      -- 
    ra_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_0, ack => convTranspose_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_320_Update/ca
      -- 
    ca_690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_1, ack => convTranspose_CP_0_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_update_start_
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Update/cr
      -- 
    ra_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_328_inst_ack_0, ack => convTranspose_CP_0_elements(94)); -- 
    cr_703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(94), ack => RPIPE_ConvTranspose_input_pipe_328_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_328_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Sample/rr
      -- 
    ca_704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_328_inst_ack_1, ack => convTranspose_CP_0_elements(95)); -- 
    rr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(95), ack => type_cast_332_inst_req_0); -- 
    rr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(95), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Sample/ra
      -- 
    ra_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_0, ack => convTranspose_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_332_Update/ca
      -- 
    ca_718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_1, ack => convTranspose_CP_0_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_update_start_
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Update/cr
      -- 
    ra_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_0, ack => convTranspose_CP_0_elements(98)); -- 
    cr_731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(98), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_341_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Sample/rr
      -- 
    ca_732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_1, ack => convTranspose_CP_0_elements(99)); -- 
    rr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(99), ack => type_cast_345_inst_req_0); -- 
    rr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(99), ack => RPIPE_ConvTranspose_input_pipe_353_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Sample/ra
      -- 
    ra_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => convTranspose_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_345_Update/ca
      -- 
    ca_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => convTranspose_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_update_start_
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Update/cr
      -- 
    ra_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_353_inst_ack_0, ack => convTranspose_CP_0_elements(102)); -- 
    cr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(102), ack => RPIPE_ConvTranspose_input_pipe_353_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_353_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Sample/$entry
      -- 
    ca_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_353_inst_ack_1, ack => convTranspose_CP_0_elements(103)); -- 
    rr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(103), ack => type_cast_357_inst_req_0); -- 
    rr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(103), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Sample/$exit
      -- 
    ra_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => convTranspose_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_357_update_completed_
      -- 
    ca_774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => convTranspose_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_update_start_
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Update/cr
      -- 
    ra_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_0, ack => convTranspose_CP_0_elements(106)); -- 
    cr_787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(106), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_366_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Sample/rr
      -- 
    ca_788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_1, ack => convTranspose_CP_0_elements(107)); -- 
    rr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(107), ack => type_cast_370_inst_req_0); -- 
    rr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(107), ack => RPIPE_ConvTranspose_input_pipe_378_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Sample/ra
      -- 
    ra_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => convTranspose_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_370_Update/ca
      -- 
    ca_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => convTranspose_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_update_start_
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Update/cr
      -- 
    ra_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_378_inst_ack_0, ack => convTranspose_CP_0_elements(110)); -- 
    cr_815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(110), ack => RPIPE_ConvTranspose_input_pipe_378_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_378_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Sample/rr
      -- 
    ca_816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_378_inst_ack_1, ack => convTranspose_CP_0_elements(111)); -- 
    rr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(111), ack => type_cast_382_inst_req_0); -- 
    rr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(111), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Sample/ra
      -- 
    ra_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_382_inst_ack_0, ack => convTranspose_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_382_Update/ca
      -- 
    ca_830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_382_inst_ack_1, ack => convTranspose_CP_0_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_update_start_
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Update/cr
      -- 
    ra_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_0, ack => convTranspose_CP_0_elements(114)); -- 
    cr_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(114), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/RPIPE_ConvTranspose_input_pipe_391_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Sample/rr
      -- 
    ca_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_1, ack => convTranspose_CP_0_elements(115)); -- 
    rr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(115), ack => type_cast_395_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Sample/ra
      -- 
    ra_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_0, ack => convTranspose_CP_0_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/type_cast_395_Update/ca
      -- 
    ca_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_1, ack => convTranspose_CP_0_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408__exit__
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_409__entry__
      -- CP-element group 118: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_408/$exit
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_409_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_409_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_409_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_409_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_25/R_cmp441_410_place
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_409_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_409_else_link/$entry
      -- 
    branch_req_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(118), ack => if_stmt_409_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(74) & convTranspose_CP_0_elements(77) & convTranspose_CP_0_elements(81) & convTranspose_CP_0_elements(85) & convTranspose_CP_0_elements(89) & convTranspose_CP_0_elements(93) & convTranspose_CP_0_elements(97) & convTranspose_CP_0_elements(68) & convTranspose_CP_0_elements(65) & convTranspose_CP_0_elements(71) & convTranspose_CP_0_elements(62) & convTranspose_CP_0_elements(59) & convTranspose_CP_0_elements(101) & convTranspose_CP_0_elements(105) & convTranspose_CP_0_elements(109) & convTranspose_CP_0_elements(113) & convTranspose_CP_0_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_430__exit__
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459__entry__
      -- CP-element group 119: 	 branch_block_stmt_25/if_stmt_409_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_25/if_stmt_409_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_25/entry_bbx_xnph443
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_update_start_
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_430_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_25/entry_bbx_xnph443_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/entry_bbx_xnph443_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_430_PhiAck/dummy
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_430_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_430_PhiAck/$entry
      -- 
    if_choice_transition_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_409_branch_ack_1, ack => convTranspose_CP_0_elements(119)); -- 
    rr_910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(119), ack => type_cast_445_inst_req_0); -- 
    cr_915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(119), ack => type_cast_445_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	430 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_25/if_stmt_409_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_25/if_stmt_409_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_25/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_25/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_25/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_409_branch_ack_0, ack => convTranspose_CP_0_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	430 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_25/merge_stmt_631_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_25/merge_stmt_631__exit__
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666__entry__
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_update_start_
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/$entry
      -- CP-element group 121: 	 branch_block_stmt_25/if_stmt_424_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_25/if_stmt_424_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_25/forx_xcond190x_xpreheader_bbx_xnph439
      -- CP-element group 121: 	 branch_block_stmt_25/merge_stmt_631_PhiAck/dummy
      -- CP-element group 121: 	 branch_block_stmt_25/merge_stmt_631_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_25/merge_stmt_631_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_25/forx_xcond190x_xpreheader_bbx_xnph439_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_25/forx_xcond190x_xpreheader_bbx_xnph439_PhiReq/$entry
      -- 
    if_choice_transition_893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_424_branch_ack_1, ack => convTranspose_CP_0_elements(121)); -- 
    cr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(121), ack => type_cast_652_inst_req_1); -- 
    rr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(121), ack => type_cast_652_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	430 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	443 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_25/if_stmt_424_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_25/if_stmt_424_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_25/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_25/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_25/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_424_branch_ack_0, ack => convTranspose_CP_0_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Sample/ra
      -- 
    ra_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_445_inst_ack_0, ack => convTranspose_CP_0_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	431 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459__exit__
      -- CP-element group 124: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/$exit
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_436_to_assign_stmt_459/type_cast_445_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/phi_stmt_462/$entry
      -- CP-element group 124: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/$entry
      -- 
    ca_916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_445_inst_ack_1, ack => convTranspose_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	436 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Sample/ack
      -- 
    ack_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_474_index_offset_ack_0, ack => convTranspose_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	436 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_request/req
      -- 
    ack_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_474_index_offset_ack_1, ack => convTranspose_CP_0_elements(126)); -- 
    req_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(126), ack => addr_of_475_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_request/ack
      -- 
    ack_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_475_final_reg_ack_0, ack => convTranspose_CP_0_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	436 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_complete/ack
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_update_completed_
      -- 
    ack_965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_475_final_reg_ack_1, ack => convTranspose_CP_0_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	436 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_update_start_
      -- 
    ra_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_478_inst_ack_0, ack => convTranspose_CP_0_elements(129)); -- 
    cr_978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(129), ack => RPIPE_ConvTranspose_input_pipe_478_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_update_completed_
      -- 
    ca_979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_478_inst_ack_1, ack => convTranspose_CP_0_elements(130)); -- 
    rr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(130), ack => type_cast_482_inst_req_0); -- 
    rr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(130), ack => RPIPE_ConvTranspose_input_pipe_491_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Sample/$exit
      -- 
    ra_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_482_inst_ack_0, ack => convTranspose_CP_0_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	436 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Update/$exit
      -- 
    ca_993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_482_inst_ack_1, ack => convTranspose_CP_0_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_update_start_
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_sample_completed_
      -- 
    ra_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_491_inst_ack_0, ack => convTranspose_CP_0_elements(133)); -- 
    cr_1006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(133), ack => RPIPE_ConvTranspose_input_pipe_491_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_491_update_completed_
      -- 
    ca_1007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_491_inst_ack_1, ack => convTranspose_CP_0_elements(134)); -- 
    rr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(134), ack => type_cast_495_inst_req_0); -- 
    rr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(134), ack => RPIPE_ConvTranspose_input_pipe_509_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_sample_completed_
      -- 
    ra_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_495_inst_ack_0, ack => convTranspose_CP_0_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	436 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_update_completed_
      -- 
    ca_1021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_495_inst_ack_1, ack => convTranspose_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_update_start_
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_sample_completed_
      -- 
    ra_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_509_inst_ack_0, ack => convTranspose_CP_0_elements(137)); -- 
    cr_1034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(137), ack => RPIPE_ConvTranspose_input_pipe_509_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_509_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Sample/$entry
      -- 
    ca_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_509_inst_ack_1, ack => convTranspose_CP_0_elements(138)); -- 
    rr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(138), ack => type_cast_513_inst_req_0); -- 
    rr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(138), ack => RPIPE_ConvTranspose_input_pipe_527_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Sample/$exit
      -- 
    ra_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_513_inst_ack_0, ack => convTranspose_CP_0_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	436 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_update_completed_
      -- 
    ca_1049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_513_inst_ack_1, ack => convTranspose_CP_0_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_update_start_
      -- 
    ra_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_527_inst_ack_0, ack => convTranspose_CP_0_elements(141)); -- 
    cr_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(141), ack => RPIPE_ConvTranspose_input_pipe_527_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_527_update_completed_
      -- 
    ca_1063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_527_inst_ack_1, ack => convTranspose_CP_0_elements(142)); -- 
    rr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(142), ack => type_cast_531_inst_req_0); -- 
    rr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(142), ack => RPIPE_ConvTranspose_input_pipe_545_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_sample_completed_
      -- 
    ra_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_0, ack => convTranspose_CP_0_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	436 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_update_completed_
      -- 
    ca_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_1, ack => convTranspose_CP_0_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_update_start_
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Sample/$exit
      -- 
    ra_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_545_inst_ack_0, ack => convTranspose_CP_0_elements(145)); -- 
    cr_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(145), ack => RPIPE_ConvTranspose_input_pipe_545_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_545_Update/$exit
      -- 
    ca_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_545_inst_ack_1, ack => convTranspose_CP_0_elements(146)); -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(146), ack => type_cast_549_inst_req_0); -- 
    rr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(146), ack => RPIPE_ConvTranspose_input_pipe_563_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_sample_completed_
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_549_inst_ack_0, ack => convTranspose_CP_0_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	436 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_update_completed_
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_549_inst_ack_1, ack => convTranspose_CP_0_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_update_start_
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_sample_completed_
      -- 
    ra_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_563_inst_ack_0, ack => convTranspose_CP_0_elements(149)); -- 
    cr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(149), ack => RPIPE_ConvTranspose_input_pipe_563_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_563_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_sample_start_
      -- 
    ca_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_563_inst_ack_1, ack => convTranspose_CP_0_elements(150)); -- 
    rr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(150), ack => type_cast_567_inst_req_0); -- 
    rr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(150), ack => RPIPE_ConvTranspose_input_pipe_581_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_sample_completed_
      -- 
    ra_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_567_inst_ack_0, ack => convTranspose_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	436 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Update/ca
      -- 
    ca_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_567_inst_ack_1, ack => convTranspose_CP_0_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_update_start_
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_sample_completed_
      -- 
    ra_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_581_inst_ack_0, ack => convTranspose_CP_0_elements(153)); -- 
    cr_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(153), ack => RPIPE_ConvTranspose_input_pipe_581_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_581_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Sample/rr
      -- 
    ca_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_581_inst_ack_1, ack => convTranspose_CP_0_elements(154)); -- 
    rr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(154), ack => type_cast_585_inst_req_0); -- 
    rr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(154), ack => RPIPE_ConvTranspose_input_pipe_599_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_sample_completed_
      -- 
    ra_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_0, ack => convTranspose_CP_0_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	436 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_update_completed_
      -- 
    ca_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_1, ack => convTranspose_CP_0_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_update_start_
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Sample/$exit
      -- 
    ra_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_599_inst_ack_0, ack => convTranspose_CP_0_elements(157)); -- 
    cr_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(157), ack => RPIPE_ConvTranspose_input_pipe_599_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_599_Update/ca
      -- 
    ca_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_599_inst_ack_1, ack => convTranspose_CP_0_elements(158)); -- 
    rr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(158), ack => type_cast_603_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_sample_completed_
      -- 
    ra_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_603_inst_ack_0, ack => convTranspose_CP_0_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	436 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_update_completed_
      -- 
    ca_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_603_inst_ack_1, ack => convTranspose_CP_0_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/ptr_deref_611_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/ptr_deref_611_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/ptr_deref_611_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/ptr_deref_611_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/$entry
      -- 
    rr_1227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(161), ack => ptr_deref_611_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(128) & convTranspose_CP_0_elements(132) & convTranspose_CP_0_elements(136) & convTranspose_CP_0_elements(140) & convTranspose_CP_0_elements(144) & convTranspose_CP_0_elements(148) & convTranspose_CP_0_elements(152) & convTranspose_CP_0_elements(156) & convTranspose_CP_0_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Sample/$exit
      -- 
    ra_1228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_611_store_0_ack_0, ack => convTranspose_CP_0_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	436 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/$exit
      -- 
    ca_1239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_611_store_0_ack_1, ack => convTranspose_CP_0_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	125 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624__exit__
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_625__entry__
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_625_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_625_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/R_exitcond3_626_place
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_625_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_625_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_625_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_625_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/$exit
      -- 
    branch_req_1247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(164), ack => if_stmt_625_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(125) & convTranspose_CP_0_elements(163);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	430 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_25/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_25/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_25/merge_stmt_415__exit__
      -- CP-element group 165: 	 branch_block_stmt_25/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_25/if_stmt_625_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_25/if_stmt_625_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_25/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_25/merge_stmt_415_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_25/merge_stmt_415_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_25/merge_stmt_415_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_25/merge_stmt_415_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_25/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_25/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_625_branch_ack_1, ack => convTranspose_CP_0_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	432 
    -- CP-element group 166: 	433 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_25/if_stmt_625_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_25/if_stmt_625_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Update/cr
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_625_branch_ack_0, ack => convTranspose_CP_0_elements(166)); -- 
    cr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(166), ack => type_cast_468_inst_req_1); -- 
    rr_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(166), ack => type_cast_468_inst_req_0); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_sample_completed_
      -- 
    ra_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_0, ack => convTranspose_CP_0_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	437 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666__exit__
      -- CP-element group 168: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/$exit
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/$entry
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_637_to_assign_stmt_666/type_cast_652_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/phi_stmt_669/$entry
      -- CP-element group 168: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/$entry
      -- 
    ca_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_1, ack => convTranspose_CP_0_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	442 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_sample_complete
      -- 
    ack_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_681_index_offset_ack_0, ack => convTranspose_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	442 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_request/req
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Update/$exit
      -- 
    ack_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_681_index_offset_ack_1, ack => convTranspose_CP_0_elements(170)); -- 
    req_1318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(170), ack => addr_of_682_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_request/ack
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_request/$exit
      -- 
    ack_1319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_682_final_reg_ack_0, ack => convTranspose_CP_0_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	442 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_word_addrgen/root_register_ack
      -- 
    ack_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_682_final_reg_ack_1, ack => convTranspose_CP_0_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	442 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_update_start_
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Update/cr
      -- 
    ra_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_685_inst_ack_0, ack => convTranspose_CP_0_elements(173)); -- 
    cr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(173), ack => RPIPE_ConvTranspose_input_pipe_685_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Update/$exit
      -- 
    ca_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_685_inst_ack_1, ack => convTranspose_CP_0_elements(174)); -- 
    rr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(174), ack => type_cast_689_inst_req_0); -- 
    rr_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(174), ack => RPIPE_ConvTranspose_input_pipe_698_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Sample/ra
      -- 
    ra_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_0, ack => convTranspose_CP_0_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	442 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Update/$exit
      -- 
    ca_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_1, ack => convTranspose_CP_0_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_update_start_
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_sample_completed_
      -- 
    ra_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_698_inst_ack_0, ack => convTranspose_CP_0_elements(177)); -- 
    cr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(177), ack => RPIPE_ConvTranspose_input_pipe_698_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_698_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_sample_start_
      -- 
    ca_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_698_inst_ack_1, ack => convTranspose_CP_0_elements(178)); -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(178), ack => type_cast_702_inst_req_0); -- 
    rr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(178), ack => RPIPE_ConvTranspose_input_pipe_716_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Sample/$exit
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_702_inst_ack_0, ack => convTranspose_CP_0_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	442 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_update_completed_
      -- 
    ca_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_702_inst_ack_1, ack => convTranspose_CP_0_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_update_start_
      -- 
    ra_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_716_inst_ack_0, ack => convTranspose_CP_0_elements(181)); -- 
    cr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(181), ack => RPIPE_ConvTranspose_input_pipe_716_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_716_Update/$exit
      -- 
    ca_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_716_inst_ack_1, ack => convTranspose_CP_0_elements(182)); -- 
    rr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(182), ack => type_cast_720_inst_req_0); -- 
    rr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(182), ack => RPIPE_ConvTranspose_input_pipe_734_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_sample_completed_
      -- 
    ra_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_720_inst_ack_0, ack => convTranspose_CP_0_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	442 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_update_completed_
      -- 
    ca_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_720_inst_ack_1, ack => convTranspose_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_update_start_
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Sample/$exit
      -- 
    ra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_734_inst_ack_0, ack => convTranspose_CP_0_elements(185)); -- 
    cr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(185), ack => RPIPE_ConvTranspose_input_pipe_734_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_734_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Sample/rr
      -- 
    ca_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_734_inst_ack_1, ack => convTranspose_CP_0_elements(186)); -- 
    rr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(186), ack => type_cast_738_inst_req_0); -- 
    rr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(186), ack => RPIPE_ConvTranspose_input_pipe_752_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Sample/ra
      -- 
    ra_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_738_inst_ack_0, ack => convTranspose_CP_0_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	442 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Update/ca
      -- 
    ca_1436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_738_inst_ack_1, ack => convTranspose_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_update_start_
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Update/cr
      -- 
    ra_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_752_inst_ack_0, ack => convTranspose_CP_0_elements(189)); -- 
    cr_1449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(189), ack => RPIPE_ConvTranspose_input_pipe_752_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_752_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Sample/rr
      -- 
    ca_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_752_inst_ack_1, ack => convTranspose_CP_0_elements(190)); -- 
    rr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(190), ack => type_cast_756_inst_req_0); -- 
    rr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(190), ack => RPIPE_ConvTranspose_input_pipe_770_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Sample/ra
      -- 
    ra_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_756_inst_ack_0, ack => convTranspose_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	442 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Update/ca
      -- 
    ca_1464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_756_inst_ack_1, ack => convTranspose_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_update_start_
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Update/cr
      -- 
    ra_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_770_inst_ack_0, ack => convTranspose_CP_0_elements(193)); -- 
    cr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(193), ack => RPIPE_ConvTranspose_input_pipe_770_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_770_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Sample/rr
      -- 
    ca_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_770_inst_ack_1, ack => convTranspose_CP_0_elements(194)); -- 
    rr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(194), ack => type_cast_774_inst_req_0); -- 
    rr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(194), ack => RPIPE_ConvTranspose_input_pipe_788_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Sample/ra
      -- 
    ra_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_774_inst_ack_0, ack => convTranspose_CP_0_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	442 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Update/ca
      -- 
    ca_1492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_774_inst_ack_1, ack => convTranspose_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_update_start_
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Update/cr
      -- 
    ra_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_788_inst_ack_0, ack => convTranspose_CP_0_elements(197)); -- 
    cr_1505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(197), ack => RPIPE_ConvTranspose_input_pipe_788_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_788_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Sample/rr
      -- 
    ca_1506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_788_inst_ack_1, ack => convTranspose_CP_0_elements(198)); -- 
    rr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(198), ack => type_cast_792_inst_req_0); -- 
    rr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(198), ack => RPIPE_ConvTranspose_input_pipe_806_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Sample/ra
      -- 
    ra_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_792_inst_ack_0, ack => convTranspose_CP_0_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	442 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Update/ca
      -- 
    ca_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_792_inst_ack_1, ack => convTranspose_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_update_start_
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Update/cr
      -- 
    ra_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_806_inst_ack_0, ack => convTranspose_CP_0_elements(201)); -- 
    cr_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(201), ack => RPIPE_ConvTranspose_input_pipe_806_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_806_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Sample/rr
      -- 
    ca_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_806_inst_ack_1, ack => convTranspose_CP_0_elements(202)); -- 
    rr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(202), ack => type_cast_810_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Sample/ra
      -- 
    ra_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_810_inst_ack_0, ack => convTranspose_CP_0_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	442 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Update/ca
      -- 
    ca_1548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_810_inst_ack_1, ack => convTranspose_CP_0_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/ptr_deref_818_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/ptr_deref_818_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/ptr_deref_818_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/ptr_deref_818_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/word_access_start/word_0/rr
      -- 
    rr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(205), ack => ptr_deref_818_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(172) & convTranspose_CP_0_elements(176) & convTranspose_CP_0_elements(180) & convTranspose_CP_0_elements(184) & convTranspose_CP_0_elements(188) & convTranspose_CP_0_elements(192) & convTranspose_CP_0_elements(196) & convTranspose_CP_0_elements(200) & convTranspose_CP_0_elements(204);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Sample/word_access_start/word_0/ra
      -- 
    ra_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_818_store_0_ack_0, ack => convTranspose_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	442 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/word_access_complete/word_0/ca
      -- 
    ca_1598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_818_store_0_ack_1, ack => convTranspose_CP_0_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	169 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831__exit__
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_832__entry__
      -- CP-element group 208: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/$exit
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_832_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_832_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_832_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_832_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_25/R_exitcond2_833_place
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_832_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_832_else_link/$entry
      -- 
    branch_req_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(208), ack => if_stmt_832_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(169) & convTranspose_CP_0_elements(207);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	443 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_838__exit__
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_838_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_838_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_838_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_25/if_stmt_832_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_25/if_stmt_832_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_838_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- 
    if_choice_transition_1611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_832_branch_ack_1, ack => convTranspose_CP_0_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	438 
    -- CP-element group 210: 	439 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/$entry
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/$entry
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_25/if_stmt_832_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_25/if_stmt_832_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_832_branch_ack_0, ack => convTranspose_CP_0_elements(210)); -- 
    cr_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(210), ack => type_cast_672_inst_req_1); -- 
    rr_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(210), ack => type_cast_672_inst_req_0); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	443 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Sample/ra
      -- 
    ra_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_0, ack => convTranspose_CP_0_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	443 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Update/ca
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_1, ack => convTranspose_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	443 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Sample/ra
      -- 
    ra_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_0, ack => convTranspose_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	443 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Update/ca
      -- 
    ca_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_1, ack => convTranspose_CP_0_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	443 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Sample/ra
      -- 
    ra_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => convTranspose_CP_0_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	443 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Update/ca
      -- 
    ca_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => convTranspose_CP_0_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868__exit__
      -- CP-element group 217: 	 branch_block_stmt_25/if_stmt_869__entry__
      -- CP-element group 217: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/$exit
      -- CP-element group 217: 	 branch_block_stmt_25/if_stmt_869_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_25/if_stmt_869_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_25/if_stmt_869_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_25/if_stmt_869_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_25/R_cmp264433_870_place
      -- CP-element group 217: 	 branch_block_stmt_25/if_stmt_869_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_25/if_stmt_869_else_link/$entry
      -- 
    branch_req_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(217), ack => if_stmt_869_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(212) & convTranspose_CP_0_elements(214) & convTranspose_CP_0_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_25/merge_stmt_875_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_25/merge_stmt_875__exit__
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910__entry__
      -- CP-element group 218: 	 branch_block_stmt_25/if_stmt_869_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_25/if_stmt_869_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_25/forx_xend250_bbx_xnph435
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/$entry
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_update_start_
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_25/merge_stmt_875_PhiAck/dummy
      -- CP-element group 218: 	 branch_block_stmt_25/merge_stmt_875_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_25/merge_stmt_875_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_25/forx_xend250_bbx_xnph435_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_25/forx_xend250_bbx_xnph435_PhiReq/$entry
      -- 
    if_choice_transition_1675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_869_branch_ack_1, ack => convTranspose_CP_0_elements(218)); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(218), ack => type_cast_896_inst_req_0); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(218), ack => type_cast_896_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	450 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_869_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_869_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_25/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_25/forx_xend250_forx_xend273_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_25/forx_xend250_forx_xend273_PhiReq/$entry
      -- 
    else_choice_transition_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_869_branch_ack_0, ack => convTranspose_CP_0_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_0, ack => convTranspose_CP_0_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	444 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910__exit__
      -- CP-element group 221: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/$exit
      -- CP-element group 221: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_25/assign_stmt_881_to_assign_stmt_910/type_cast_896_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/phi_stmt_913/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/$entry
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_1, ack => convTranspose_CP_0_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	449 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Sample/ack
      -- 
    ack_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_925_index_offset_ack_0, ack => convTranspose_CP_0_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	449 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_request/req
      -- 
    ack_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_925_index_offset_ack_1, ack => convTranspose_CP_0_elements(223)); -- 
    req_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(223), ack => addr_of_926_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_request/ack
      -- 
    ack_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_926_final_reg_ack_0, ack => convTranspose_CP_0_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	449 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/ptr_deref_929_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/ptr_deref_929_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/ptr_deref_929_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/ptr_deref_929_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/word_access_start/word_0/rr
      -- 
    ack_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_926_final_reg_ack_1, ack => convTranspose_CP_0_elements(225)); -- 
    rr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(225), ack => ptr_deref_929_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Sample/word_access_start/word_0/ra
      -- 
    ra_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_929_store_0_ack_0, ack => convTranspose_CP_0_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	449 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/word_access_complete/word_0/ca
      -- 
    ca_1797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_929_store_0_ack_1, ack => convTranspose_CP_0_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943__exit__
      -- CP-element group 228: 	 branch_block_stmt_25/if_stmt_944__entry__
      -- CP-element group 228: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/$exit
      -- CP-element group 228: 	 branch_block_stmt_25/if_stmt_944_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_25/if_stmt_944_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_25/if_stmt_944_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_25/if_stmt_944_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_25/R_exitcond_945_place
      -- CP-element group 228: 	 branch_block_stmt_25/if_stmt_944_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_25/if_stmt_944_else_link/$entry
      -- 
    branch_req_1805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(228), ack => if_stmt_944_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(222) & convTranspose_CP_0_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	450 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_25/merge_stmt_950__exit__
      -- CP-element group 229: 	 branch_block_stmt_25/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_25/merge_stmt_950_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_25/if_stmt_944_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_25/if_stmt_944_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_25/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_25/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_25/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_25/merge_stmt_950_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_25/merge_stmt_950_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_25/merge_stmt_950_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_25/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_25/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_944_branch_ack_1, ack => convTranspose_CP_0_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	445 
    -- CP-element group 230: 	446 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_25/if_stmt_944_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_25/if_stmt_944_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/$entry
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/$entry
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_944_branch_ack_0, ack => convTranspose_CP_0_elements(230)); -- 
    rr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(230), ack => type_cast_916_inst_req_0); -- 
    cr_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(230), ack => type_cast_916_inst_req_1); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	450 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (6) 
      -- CP-element group 231: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_update_start_
      -- CP-element group 231: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Sample/ack
      -- CP-element group 231: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Update/req
      -- 
    ack_1828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_954_inst_ack_0, ack => convTranspose_CP_0_elements(231)); -- 
    req_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(231), ack => WPIPE_ConvTranspose_output_pipe_954_inst_req_1); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Update/ack
      -- CP-element group 232: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Sample/req
      -- 
    ack_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_954_inst_ack_1, ack => convTranspose_CP_0_elements(232)); -- 
    req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(232), ack => WPIPE_ConvTranspose_output_pipe_958_inst_req_0); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_update_start_
      -- CP-element group 233: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Sample/ack
      -- CP-element group 233: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Update/req
      -- 
    ack_1842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_958_inst_ack_0, ack => convTranspose_CP_0_elements(233)); -- 
    req_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(233), ack => WPIPE_ConvTranspose_output_pipe_958_inst_req_1); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	263 
    -- CP-element group 234: 	281 
    -- CP-element group 234: 	282 
    -- CP-element group 234: 	286 
    -- CP-element group 234: 	287 
    -- CP-element group 234: 	297 
    -- CP-element group 234: 	315 
    -- CP-element group 234: 	316 
    -- CP-element group 234: 	320 
    -- CP-element group 234: 	321 
    -- CP-element group 234: 	331 
    -- CP-element group 234: 	349 
    -- CP-element group 234: 	350 
    -- CP-element group 234: 	354 
    -- CP-element group 234: 	355 
    -- CP-element group 234: 	365 
    -- CP-element group 234: 	367 
    -- CP-element group 234: 	369 
    -- CP-element group 234: 	371 
    -- CP-element group 234:  members (67) 
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961__exit__
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186__entry__
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_update_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_update_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_update_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_update_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/$exit
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_958_Update/ack
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_update_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_update_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Sample/rr
      -- 
    ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_958_inst_ack_1, ack => convTranspose_CP_0_elements(234)); -- 
    cr_2213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1049_inst_req_1); -- 
    cr_2185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1042_inst_req_1); -- 
    req_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => WPIPE_Block1_start_1007_inst_req_0); -- 
    rr_2208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1049_inst_req_0); -- 
    cr_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1098_inst_req_1); -- 
    rr_2180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1042_inst_req_0); -- 
    rr_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1098_inst_req_0); -- 
    cr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1105_inst_req_1); -- 
    req_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => WPIPE_Block2_start_1063_inst_req_0); -- 
    rr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1105_inst_req_0); -- 
    req_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => WPIPE_Block0_start_963_inst_req_0); -- 
    req_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => WPIPE_Block3_start_1119_inst_req_0); -- 
    rr_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1154_inst_req_0); -- 
    cr_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1154_inst_req_1); -- 
    rr_2656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1161_inst_req_0); -- 
    cr_2661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => type_cast_1161_inst_req_1); -- 
    rr_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => RPIPE_Block0_done_1176_inst_req_0); -- 
    rr_2740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => RPIPE_Block1_done_1179_inst_req_0); -- 
    rr_2754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => RPIPE_Block2_done_1182_inst_req_0); -- 
    rr_2768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(234), ack => RPIPE_Block3_done_1185_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_update_start_
      -- CP-element group 235: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Update/req
      -- 
    ack_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_963_inst_ack_0, ack => convTranspose_CP_0_elements(235)); -- 
    req_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(235), ack => WPIPE_Block0_start_963_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_963_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Sample/req
      -- 
    ack_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_963_inst_ack_1, ack => convTranspose_CP_0_elements(236)); -- 
    req_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(236), ack => WPIPE_Block0_start_966_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_update_start_
      -- CP-element group 237: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Update/req
      -- 
    ack_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_966_inst_ack_0, ack => convTranspose_CP_0_elements(237)); -- 
    req_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(237), ack => WPIPE_Block0_start_966_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_966_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Sample/req
      -- 
    ack_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_966_inst_ack_1, ack => convTranspose_CP_0_elements(238)); -- 
    req_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(238), ack => WPIPE_Block0_start_969_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_update_start_
      -- CP-element group 239: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Update/req
      -- 
    ack_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_969_inst_ack_0, ack => convTranspose_CP_0_elements(239)); -- 
    req_1891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(239), ack => WPIPE_Block0_start_969_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_969_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Sample/req
      -- 
    ack_1892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_969_inst_ack_1, ack => convTranspose_CP_0_elements(240)); -- 
    req_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(240), ack => WPIPE_Block0_start_972_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_update_start_
      -- CP-element group 241: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Update/req
      -- 
    ack_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_972_inst_ack_0, ack => convTranspose_CP_0_elements(241)); -- 
    req_1905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(241), ack => WPIPE_Block0_start_972_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_972_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/req
      -- 
    ack_1906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_972_inst_ack_1, ack => convTranspose_CP_0_elements(242)); -- 
    req_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(242), ack => WPIPE_Block0_start_975_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_update_start_
      -- CP-element group 243: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/req
      -- 
    ack_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_0, ack => convTranspose_CP_0_elements(243)); -- 
    req_1919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(243), ack => WPIPE_Block0_start_975_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/req
      -- 
    ack_1920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_1, ack => convTranspose_CP_0_elements(244)); -- 
    req_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(244), ack => WPIPE_Block0_start_978_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_update_start_
      -- CP-element group 245: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/req
      -- 
    ack_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_0, ack => convTranspose_CP_0_elements(245)); -- 
    req_1933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(245), ack => WPIPE_Block0_start_978_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/req
      -- 
    ack_1934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_1, ack => convTranspose_CP_0_elements(246)); -- 
    req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(246), ack => WPIPE_Block0_start_981_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_update_start_
      -- CP-element group 247: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/req
      -- 
    ack_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_0, ack => convTranspose_CP_0_elements(247)); -- 
    req_1947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(247), ack => WPIPE_Block0_start_981_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/req
      -- 
    ack_1948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_1, ack => convTranspose_CP_0_elements(248)); -- 
    req_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(248), ack => WPIPE_Block0_start_984_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_update_start_
      -- CP-element group 249: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/req
      -- 
    ack_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_0, ack => convTranspose_CP_0_elements(249)); -- 
    req_1961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(249), ack => WPIPE_Block0_start_984_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/req
      -- 
    ack_1962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_1, ack => convTranspose_CP_0_elements(250)); -- 
    req_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(250), ack => WPIPE_Block0_start_987_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_update_start_
      -- CP-element group 251: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/req
      -- 
    ack_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_0, ack => convTranspose_CP_0_elements(251)); -- 
    req_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(251), ack => WPIPE_Block0_start_987_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/req
      -- 
    ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_1, ack => convTranspose_CP_0_elements(252)); -- 
    req_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(252), ack => WPIPE_Block0_start_990_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_update_start_
      -- CP-element group 253: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/req
      -- 
    ack_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_0, ack => convTranspose_CP_0_elements(253)); -- 
    req_1989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(253), ack => WPIPE_Block0_start_990_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Sample/req
      -- 
    ack_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_1, ack => convTranspose_CP_0_elements(254)); -- 
    req_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(254), ack => WPIPE_Block0_start_994_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Update/req
      -- CP-element group 255: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_update_start_
      -- CP-element group 255: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Sample/ack
      -- 
    ack_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_0, ack => convTranspose_CP_0_elements(255)); -- 
    req_2003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(255), ack => WPIPE_Block0_start_994_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_994_update_completed_
      -- 
    ack_2004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_1, ack => convTranspose_CP_0_elements(256)); -- 
    req_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(256), ack => WPIPE_Block0_start_998_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Update/req
      -- CP-element group 257: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_update_start_
      -- CP-element group 257: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_sample_completed_
      -- 
    ack_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_998_inst_ack_0, ack => convTranspose_CP_0_elements(257)); -- 
    req_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(257), ack => WPIPE_Block0_start_998_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_998_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Sample/req
      -- 
    ack_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_998_inst_ack_1, ack => convTranspose_CP_0_elements(258)); -- 
    req_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(258), ack => WPIPE_Block0_start_1001_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_update_start_
      -- CP-element group 259: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Update/req
      -- CP-element group 259: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Sample/ack
      -- 
    ack_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1001_inst_ack_0, ack => convTranspose_CP_0_elements(259)); -- 
    req_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(259), ack => WPIPE_Block0_start_1001_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1001_Update/$exit
      -- 
    ack_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1001_inst_ack_1, ack => convTranspose_CP_0_elements(260)); -- 
    req_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(260), ack => WPIPE_Block0_start_1004_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Update/req
      -- CP-element group 261: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_update_start_
      -- CP-element group 261: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_sample_completed_
      -- 
    ack_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1004_inst_ack_0, ack => convTranspose_CP_0_elements(261)); -- 
    req_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(261), ack => WPIPE_Block0_start_1004_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	373 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block0_start_1004_update_completed_
      -- 
    ack_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1004_inst_ack_1, ack => convTranspose_CP_0_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	234 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_update_start_
      -- CP-element group 263: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Update/req
      -- CP-element group 263: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Update/$entry
      -- 
    ack_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1007_inst_ack_0, ack => convTranspose_CP_0_elements(263)); -- 
    req_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(263), ack => WPIPE_Block1_start_1007_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Sample/req
      -- CP-element group 264: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1007_Update/$exit
      -- 
    ack_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1007_inst_ack_1, ack => convTranspose_CP_0_elements(264)); -- 
    req_2068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(264), ack => WPIPE_Block1_start_1010_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Update/req
      -- CP-element group 265: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_update_start_
      -- CP-element group 265: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_sample_completed_
      -- 
    ack_2069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1010_inst_ack_0, ack => convTranspose_CP_0_elements(265)); -- 
    req_2073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(265), ack => WPIPE_Block1_start_1010_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1010_update_completed_
      -- 
    ack_2074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1010_inst_ack_1, ack => convTranspose_CP_0_elements(266)); -- 
    req_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(266), ack => WPIPE_Block1_start_1013_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_update_start_
      -- CP-element group 267: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Update/req
      -- CP-element group 267: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_sample_completed_
      -- 
    ack_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_0, ack => convTranspose_CP_0_elements(267)); -- 
    req_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(267), ack => WPIPE_Block1_start_1013_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1013_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_sample_start_
      -- 
    ack_2088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_1, ack => convTranspose_CP_0_elements(268)); -- 
    req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(268), ack => WPIPE_Block1_start_1016_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_update_start_
      -- CP-element group 269: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Update/req
      -- 
    ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_0, ack => convTranspose_CP_0_elements(269)); -- 
    req_2101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(269), ack => WPIPE_Block1_start_1016_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1016_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/req
      -- 
    ack_2102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_1, ack => convTranspose_CP_0_elements(270)); -- 
    req_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(270), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_update_start_
      -- CP-element group 271: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/req
      -- CP-element group 271: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/$exit
      -- 
    ack_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_0_elements(271)); -- 
    req_2115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(271), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/$exit
      -- 
    ack_2116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_0_elements(272)); -- 
    req_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(272), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_update_start_
      -- CP-element group 273: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/req
      -- 
    ack_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_0_elements(273)); -- 
    req_2129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(273), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/ack
      -- 
    ack_2130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_0_elements(274)); -- 
    req_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(274), ack => WPIPE_Block1_start_1025_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/req
      -- CP-element group 275: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_update_start_
      -- CP-element group 275: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_sample_completed_
      -- 
    ack_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_0, ack => convTranspose_CP_0_elements(275)); -- 
    req_2143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(275), ack => WPIPE_Block1_start_1025_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1025_update_completed_
      -- 
    ack_2144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_1, ack => convTranspose_CP_0_elements(276)); -- 
    req_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(276), ack => WPIPE_Block1_start_1028_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/req
      -- CP-element group 277: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_update_start_
      -- CP-element group 277: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_sample_completed_
      -- 
    ack_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_0, ack => convTranspose_CP_0_elements(277)); -- 
    req_2157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(277), ack => WPIPE_Block1_start_1028_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1028_update_completed_
      -- 
    ack_2158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_1, ack => convTranspose_CP_0_elements(278)); -- 
    req_2166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(278), ack => WPIPE_Block1_start_1031_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/req
      -- CP-element group 279: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_update_start_
      -- CP-element group 279: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_sample_completed_
      -- 
    ack_2167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_0, ack => convTranspose_CP_0_elements(279)); -- 
    req_2171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(279), ack => WPIPE_Block1_start_1031_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1031_update_completed_
      -- 
    ack_2172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_1, ack => convTranspose_CP_0_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	234 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_sample_completed_
      -- 
    ra_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1042_inst_ack_0, ack => convTranspose_CP_0_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	234 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1042_update_completed_
      -- 
    ca_2186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1042_inst_ack_1, ack => convTranspose_CP_0_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_sample_start_
      -- 
    req_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(283), ack => WPIPE_Block1_start_1044_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(280) & convTranspose_CP_0_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Update/req
      -- CP-element group 284: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_update_start_
      -- CP-element group 284: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Sample/$exit
      -- 
    ack_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1044_inst_ack_0, ack => convTranspose_CP_0_elements(284)); -- 
    req_2199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(284), ack => WPIPE_Block1_start_1044_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_Update/ack
      -- CP-element group 285: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1044_update_completed_
      -- 
    ack_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1044_inst_ack_1, ack => convTranspose_CP_0_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	234 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Sample/ra
      -- 
    ra_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_0, ack => convTranspose_CP_0_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	234 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1049_update_completed_
      -- 
    ca_2214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_1, ack => convTranspose_CP_0_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Sample/req
      -- 
    req_2222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(288), ack => WPIPE_Block1_start_1051_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(285) & convTranspose_CP_0_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_sample_completed_
      -- CP-element group 289: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_update_start_
      -- CP-element group 289: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Update/req
      -- CP-element group 289: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Sample/ack
      -- 
    ack_2223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1051_inst_ack_0, ack => convTranspose_CP_0_elements(289)); -- 
    req_2227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(289), ack => WPIPE_Block1_start_1051_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1051_Update/$exit
      -- 
    ack_2228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1051_inst_ack_1, ack => convTranspose_CP_0_elements(290)); -- 
    req_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(290), ack => WPIPE_Block1_start_1054_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Update/req
      -- CP-element group 291: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_update_start_
      -- CP-element group 291: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_sample_completed_
      -- 
    ack_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1054_inst_ack_0, ack => convTranspose_CP_0_elements(291)); -- 
    req_2241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(291), ack => WPIPE_Block1_start_1054_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1054_update_completed_
      -- 
    ack_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1054_inst_ack_1, ack => convTranspose_CP_0_elements(292)); -- 
    req_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(292), ack => WPIPE_Block1_start_1057_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_update_start_
      -- CP-element group 293: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Update/req
      -- 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_0, ack => convTranspose_CP_0_elements(293)); -- 
    req_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(293), ack => WPIPE_Block1_start_1057_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1057_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_sample_start_
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_1, ack => convTranspose_CP_0_elements(294)); -- 
    req_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(294), ack => WPIPE_Block1_start_1060_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Update/req
      -- CP-element group 295: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_update_start_
      -- CP-element group 295: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_sample_completed_
      -- 
    ack_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1060_inst_ack_0, ack => convTranspose_CP_0_elements(295)); -- 
    req_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(295), ack => WPIPE_Block1_start_1060_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	373 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block1_start_1060_update_completed_
      -- 
    ack_2270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1060_inst_ack_1, ack => convTranspose_CP_0_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	234 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Update/req
      -- CP-element group 297: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_update_start_
      -- CP-element group 297: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_sample_completed_
      -- 
    ack_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1063_inst_ack_0, ack => convTranspose_CP_0_elements(297)); -- 
    req_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(297), ack => WPIPE_Block2_start_1063_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1063_update_completed_
      -- 
    ack_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1063_inst_ack_1, ack => convTranspose_CP_0_elements(298)); -- 
    req_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(298), ack => WPIPE_Block2_start_1066_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Update/req
      -- CP-element group 299: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_update_start_
      -- CP-element group 299: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_sample_completed_
      -- 
    ack_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1066_inst_ack_0, ack => convTranspose_CP_0_elements(299)); -- 
    req_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(299), ack => WPIPE_Block2_start_1066_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1066_update_completed_
      -- 
    ack_2298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1066_inst_ack_1, ack => convTranspose_CP_0_elements(300)); -- 
    req_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(300), ack => WPIPE_Block2_start_1069_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_update_start_
      -- CP-element group 301: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Update/req
      -- CP-element group 301: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Update/$entry
      -- 
    ack_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1069_inst_ack_0, ack => convTranspose_CP_0_elements(301)); -- 
    req_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(301), ack => WPIPE_Block2_start_1069_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1069_Update/ack
      -- 
    ack_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1069_inst_ack_1, ack => convTranspose_CP_0_elements(302)); -- 
    req_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(302), ack => WPIPE_Block2_start_1072_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Update/req
      -- CP-element group 303: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_update_start_
      -- CP-element group 303: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_sample_completed_
      -- 
    ack_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1072_inst_ack_0, ack => convTranspose_CP_0_elements(303)); -- 
    req_2325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(303), ack => WPIPE_Block2_start_1072_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1072_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_sample_start_
      -- 
    ack_2326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1072_inst_ack_1, ack => convTranspose_CP_0_elements(304)); -- 
    req_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(304), ack => WPIPE_Block2_start_1075_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/req
      -- CP-element group 305: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_update_start_
      -- CP-element group 305: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_sample_completed_
      -- 
    ack_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_0, ack => convTranspose_CP_0_elements(305)); -- 
    req_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(305), ack => WPIPE_Block2_start_1075_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1075_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/$entry
      -- 
    ack_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_1, ack => convTranspose_CP_0_elements(306)); -- 
    req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(306), ack => WPIPE_Block2_start_1078_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_update_start_
      -- CP-element group 307: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/req
      -- CP-element group 307: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/$exit
      -- 
    ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_0, ack => convTranspose_CP_0_elements(307)); -- 
    req_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(307), ack => WPIPE_Block2_start_1078_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/$exit
      -- 
    ack_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_1, ack => convTranspose_CP_0_elements(308)); -- 
    req_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(308), ack => WPIPE_Block2_start_1081_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/req
      -- CP-element group 309: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_update_start_
      -- CP-element group 309: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_sample_completed_
      -- 
    ack_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_0, ack => convTranspose_CP_0_elements(309)); -- 
    req_2367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(309), ack => WPIPE_Block2_start_1081_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1081_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_sample_start_
      -- 
    ack_2368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_1, ack => convTranspose_CP_0_elements(310)); -- 
    req_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(310), ack => WPIPE_Block2_start_1084_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/req
      -- CP-element group 311: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_update_start_
      -- CP-element group 311: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_sample_completed_
      -- 
    ack_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_0, ack => convTranspose_CP_0_elements(311)); -- 
    req_2381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(311), ack => WPIPE_Block2_start_1084_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/req
      -- CP-element group 312: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1084_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_sample_start_
      -- 
    ack_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_1, ack => convTranspose_CP_0_elements(312)); -- 
    req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(312), ack => WPIPE_Block2_start_1087_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_update_start_
      -- CP-element group 313: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/req
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_0, ack => convTranspose_CP_0_elements(313)); -- 
    req_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(313), ack => WPIPE_Block2_start_1087_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/$exit
      -- 
    ack_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_1, ack => convTranspose_CP_0_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	234 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Sample/ra
      -- CP-element group 315: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Sample/$exit
      -- 
    ra_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_0, ack => convTranspose_CP_0_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	234 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Update/ca
      -- CP-element group 316: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1098_update_completed_
      -- 
    ca_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_1, ack => convTranspose_CP_0_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Sample/req
      -- 
    req_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(317), ack => WPIPE_Block2_start_1100_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(314) & convTranspose_CP_0_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_update_start_
      -- CP-element group 318: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Update/req
      -- CP-element group 318: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Sample/ack
      -- 
    ack_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1100_inst_ack_0, ack => convTranspose_CP_0_elements(318)); -- 
    req_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(318), ack => WPIPE_Block2_start_1100_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Update/ack
      -- CP-element group 319: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1100_Update/$exit
      -- 
    ack_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1100_inst_ack_1, ack => convTranspose_CP_0_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	234 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Sample/ra
      -- CP-element group 320: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_sample_completed_
      -- 
    ra_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_0, ack => convTranspose_CP_0_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	234 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1105_Update/ca
      -- 
    ca_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_1, ack => convTranspose_CP_0_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Sample/req
      -- 
    req_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(322), ack => WPIPE_Block2_start_1107_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(319) & convTranspose_CP_0_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_update_start_
      -- CP-element group 323: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Update/req
      -- 
    ack_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1107_inst_ack_0, ack => convTranspose_CP_0_elements(323)); -- 
    req_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(323), ack => WPIPE_Block2_start_1107_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1107_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Sample/req
      -- 
    ack_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1107_inst_ack_1, ack => convTranspose_CP_0_elements(324)); -- 
    req_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(324), ack => WPIPE_Block2_start_1110_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_update_start_
      -- CP-element group 325: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Update/req
      -- 
    ack_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1110_inst_ack_0, ack => convTranspose_CP_0_elements(325)); -- 
    req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(325), ack => WPIPE_Block2_start_1110_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1110_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Sample/req
      -- 
    ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1110_inst_ack_1, ack => convTranspose_CP_0_elements(326)); -- 
    req_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(326), ack => WPIPE_Block2_start_1113_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_update_start_
      -- CP-element group 327: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Update/req
      -- 
    ack_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_0, ack => convTranspose_CP_0_elements(327)); -- 
    req_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(327), ack => WPIPE_Block2_start_1113_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1113_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Sample/req
      -- 
    ack_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_1, ack => convTranspose_CP_0_elements(328)); -- 
    req_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(328), ack => WPIPE_Block2_start_1116_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_update_start_
      -- CP-element group 329: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Update/req
      -- 
    ack_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_0, ack => convTranspose_CP_0_elements(329)); -- 
    req_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(329), ack => WPIPE_Block2_start_1116_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	373 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block2_start_1116_Update/ack
      -- 
    ack_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_1, ack => convTranspose_CP_0_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	234 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_update_start_
      -- CP-element group 331: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Update/req
      -- 
    ack_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1119_inst_ack_0, ack => convTranspose_CP_0_elements(331)); -- 
    req_2507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(331), ack => WPIPE_Block3_start_1119_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1119_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Sample/req
      -- 
    ack_2508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1119_inst_ack_1, ack => convTranspose_CP_0_elements(332)); -- 
    req_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(332), ack => WPIPE_Block3_start_1122_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_update_start_
      -- CP-element group 333: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Update/req
      -- 
    ack_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1122_inst_ack_0, ack => convTranspose_CP_0_elements(333)); -- 
    req_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(333), ack => WPIPE_Block3_start_1122_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1122_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Sample/req
      -- 
    ack_2522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1122_inst_ack_1, ack => convTranspose_CP_0_elements(334)); -- 
    req_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(334), ack => WPIPE_Block3_start_1125_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_update_start_
      -- CP-element group 335: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Update/req
      -- 
    ack_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1125_inst_ack_0, ack => convTranspose_CP_0_elements(335)); -- 
    req_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(335), ack => WPIPE_Block3_start_1125_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1125_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Sample/req
      -- 
    ack_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1125_inst_ack_1, ack => convTranspose_CP_0_elements(336)); -- 
    req_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(336), ack => WPIPE_Block3_start_1128_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_update_start_
      -- CP-element group 337: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Update/req
      -- 
    ack_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1128_inst_ack_0, ack => convTranspose_CP_0_elements(337)); -- 
    req_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(337), ack => WPIPE_Block3_start_1128_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1128_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/req
      -- 
    ack_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1128_inst_ack_1, ack => convTranspose_CP_0_elements(338)); -- 
    req_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(338), ack => WPIPE_Block3_start_1131_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_update_start_
      -- CP-element group 339: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/req
      -- 
    ack_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_0, ack => convTranspose_CP_0_elements(339)); -- 
    req_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(339), ack => WPIPE_Block3_start_1131_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/req
      -- 
    ack_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_1, ack => convTranspose_CP_0_elements(340)); -- 
    req_2572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(340), ack => WPIPE_Block3_start_1134_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_update_start_
      -- CP-element group 341: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/req
      -- 
    ack_2573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_0, ack => convTranspose_CP_0_elements(341)); -- 
    req_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(341), ack => WPIPE_Block3_start_1134_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/req
      -- 
    ack_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_1, ack => convTranspose_CP_0_elements(342)); -- 
    req_2586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(342), ack => WPIPE_Block3_start_1137_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_update_start_
      -- CP-element group 343: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/req
      -- 
    ack_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_0, ack => convTranspose_CP_0_elements(343)); -- 
    req_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(343), ack => WPIPE_Block3_start_1137_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/req
      -- 
    ack_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_1, ack => convTranspose_CP_0_elements(344)); -- 
    req_2600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(344), ack => WPIPE_Block3_start_1140_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_update_start_
      -- CP-element group 345: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/req
      -- 
    ack_2601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_0, ack => convTranspose_CP_0_elements(345)); -- 
    req_2605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(345), ack => WPIPE_Block3_start_1140_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/req
      -- 
    ack_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_1, ack => convTranspose_CP_0_elements(346)); -- 
    req_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(346), ack => WPIPE_Block3_start_1143_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_update_start_
      -- CP-element group 347: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/req
      -- 
    ack_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_0, ack => convTranspose_CP_0_elements(347)); -- 
    req_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(347), ack => WPIPE_Block3_start_1143_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/ack
      -- 
    ack_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_1, ack => convTranspose_CP_0_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	234 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Sample/ra
      -- 
    ra_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1154_inst_ack_0, ack => convTranspose_CP_0_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	234 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1154_Update/ca
      -- 
    ca_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1154_inst_ack_1, ack => convTranspose_CP_0_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Sample/req
      -- 
    req_2642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(351), ack => WPIPE_Block3_start_1156_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(348) & convTranspose_CP_0_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_update_start_
      -- CP-element group 352: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Update/req
      -- 
    ack_2643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1156_inst_ack_0, ack => convTranspose_CP_0_elements(352)); -- 
    req_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(352), ack => WPIPE_Block3_start_1156_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1156_Update/ack
      -- 
    ack_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1156_inst_ack_1, ack => convTranspose_CP_0_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	234 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Sample/ra
      -- 
    ra_2657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_0, ack => convTranspose_CP_0_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	234 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/type_cast_1161_Update/ca
      -- 
    ca_2662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_1, ack => convTranspose_CP_0_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Sample/req
      -- 
    req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(356), ack => WPIPE_Block3_start_1163_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(353) & convTranspose_CP_0_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_update_start_
      -- CP-element group 357: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Update/req
      -- 
    ack_2671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1163_inst_ack_0, ack => convTranspose_CP_0_elements(357)); -- 
    req_2675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(357), ack => WPIPE_Block3_start_1163_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1163_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Sample/req
      -- 
    ack_2676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1163_inst_ack_1, ack => convTranspose_CP_0_elements(358)); -- 
    req_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(358), ack => WPIPE_Block3_start_1166_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_update_start_
      -- CP-element group 359: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Update/req
      -- 
    ack_2685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1166_inst_ack_0, ack => convTranspose_CP_0_elements(359)); -- 
    req_2689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(359), ack => WPIPE_Block3_start_1166_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1166_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Sample/req
      -- 
    ack_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1166_inst_ack_1, ack => convTranspose_CP_0_elements(360)); -- 
    req_2698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(360), ack => WPIPE_Block3_start_1169_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_update_start_
      -- CP-element group 361: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Update/req
      -- 
    ack_2699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_0, ack => convTranspose_CP_0_elements(361)); -- 
    req_2703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(361), ack => WPIPE_Block3_start_1169_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1169_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Sample/req
      -- 
    ack_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_1, ack => convTranspose_CP_0_elements(362)); -- 
    req_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(362), ack => WPIPE_Block3_start_1172_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_update_start_
      -- CP-element group 363: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Update/req
      -- 
    ack_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_0, ack => convTranspose_CP_0_elements(363)); -- 
    req_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(363), ack => WPIPE_Block3_start_1172_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	373 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/WPIPE_Block3_start_1172_Update/ack
      -- 
    ack_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_1, ack => convTranspose_CP_0_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	234 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_update_start_
      -- CP-element group 365: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Update/cr
      -- 
    ra_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1176_inst_ack_0, ack => convTranspose_CP_0_elements(365)); -- 
    cr_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(365), ack => RPIPE_Block0_done_1176_inst_req_1); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	373 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block0_done_1176_Update/ca
      -- 
    ca_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1176_inst_ack_1, ack => convTranspose_CP_0_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	234 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_update_start_
      -- CP-element group 367: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Sample/ra
      -- CP-element group 367: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Update/cr
      -- 
    ra_2741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1179_inst_ack_0, ack => convTranspose_CP_0_elements(367)); -- 
    cr_2745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(367), ack => RPIPE_Block1_done_1179_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block1_done_1179_Update/ca
      -- 
    ca_2746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1179_inst_ack_1, ack => convTranspose_CP_0_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	234 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_update_start_
      -- CP-element group 369: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Update/cr
      -- 
    ra_2755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1182_inst_ack_0, ack => convTranspose_CP_0_elements(369)); -- 
    cr_2759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(369), ack => RPIPE_Block2_done_1182_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	373 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block2_done_1182_Update/ca
      -- 
    ca_2760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1182_inst_ack_1, ack => convTranspose_CP_0_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	234 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_update_start_
      -- CP-element group 371: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Update/cr
      -- 
    ra_2769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1185_inst_ack_0, ack => convTranspose_CP_0_elements(371)); -- 
    cr_2773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(371), ack => RPIPE_Block3_done_1185_inst_req_1); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/RPIPE_Block3_done_1185_Update/ca
      -- 
    ca_2774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1185_inst_ack_1, ack => convTranspose_CP_0_elements(372)); -- 
    -- CP-element group 373:  join  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	296 
    -- CP-element group 373: 	330 
    -- CP-element group 373: 	364 
    -- CP-element group 373: 	366 
    -- CP-element group 373: 	368 
    -- CP-element group 373: 	370 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (7) 
      -- CP-element group 373: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186__exit__
      -- CP-element group 373: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195__entry__
      -- CP-element group 373: 	 branch_block_stmt_25/assign_stmt_965_to_assign_stmt_1186/$exit
      -- CP-element group 373: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/$entry
      -- CP-element group 373: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Sample/req
      -- 
    req_2785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(373), ack => WPIPE_ConvTranspose_output_pipe_1188_inst_req_0); -- 
    convTranspose_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(262) & convTranspose_CP_0_elements(296) & convTranspose_CP_0_elements(330) & convTranspose_CP_0_elements(364) & convTranspose_CP_0_elements(366) & convTranspose_CP_0_elements(368) & convTranspose_CP_0_elements(370) & convTranspose_CP_0_elements(372);
      gj_convTranspose_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  transition  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (6) 
      -- CP-element group 374: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_update_start_
      -- CP-element group 374: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Sample/ack
      -- CP-element group 374: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Update/req
      -- 
    ack_2786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1188_inst_ack_0, ack => convTranspose_CP_0_elements(374)); -- 
    req_2790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(374), ack => WPIPE_ConvTranspose_output_pipe_1188_inst_req_1); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1188_Update/ack
      -- CP-element group 375: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Sample/req
      -- 
    ack_2791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1188_inst_ack_1, ack => convTranspose_CP_0_elements(375)); -- 
    req_2799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(375), ack => WPIPE_ConvTranspose_output_pipe_1192_inst_req_0); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_update_start_
      -- CP-element group 376: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Sample/ack
      -- CP-element group 376: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Update/req
      -- 
    ack_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1192_inst_ack_0, ack => convTranspose_CP_0_elements(376)); -- 
    req_2804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(376), ack => WPIPE_ConvTranspose_output_pipe_1192_inst_req_1); -- 
    -- CP-element group 377:  branch  transition  place  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (13) 
      -- CP-element group 377: 	 branch_block_stmt_25/if_stmt_1197__entry__
      -- CP-element group 377: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195__exit__
      -- CP-element group 377: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/$exit
      -- CP-element group 377: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1195/WPIPE_ConvTranspose_output_pipe_1192_Update/ack
      -- CP-element group 377: 	 branch_block_stmt_25/if_stmt_1197_dead_link/$entry
      -- CP-element group 377: 	 branch_block_stmt_25/if_stmt_1197_eval_test/$entry
      -- CP-element group 377: 	 branch_block_stmt_25/if_stmt_1197_eval_test/$exit
      -- CP-element group 377: 	 branch_block_stmt_25/if_stmt_1197_eval_test/branch_req
      -- CP-element group 377: 	 branch_block_stmt_25/R_cmp264433_1198_place
      -- CP-element group 377: 	 branch_block_stmt_25/if_stmt_1197_if_link/$entry
      -- CP-element group 377: 	 branch_block_stmt_25/if_stmt_1197_else_link/$entry
      -- 
    ack_2805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1192_inst_ack_1, ack => convTranspose_CP_0_elements(377)); -- 
    branch_req_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(377), ack => if_stmt_1197_branch_req_0); -- 
    -- CP-element group 378:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378: 	381 
    -- CP-element group 378:  members (18) 
      -- CP-element group 378: 	 branch_block_stmt_25/merge_stmt_1203__exit__
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238__entry__
      -- CP-element group 378: 	 branch_block_stmt_25/merge_stmt_1203_PhiReqMerge
      -- CP-element group 378: 	 branch_block_stmt_25/merge_stmt_1203_PhiAck/dummy
      -- CP-element group 378: 	 branch_block_stmt_25/merge_stmt_1203_PhiAck/$exit
      -- CP-element group 378: 	 branch_block_stmt_25/merge_stmt_1203_PhiAck/$entry
      -- CP-element group 378: 	 branch_block_stmt_25/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 378: 	 branch_block_stmt_25/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 378: 	 branch_block_stmt_25/if_stmt_1197_if_link/$exit
      -- CP-element group 378: 	 branch_block_stmt_25/if_stmt_1197_if_link/if_choice_transition
      -- CP-element group 378: 	 branch_block_stmt_25/forx_xend273_bbx_xnph
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/$entry
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_update_start_
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Update/cr
      -- 
    if_choice_transition_2818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1197_branch_ack_1, ack => convTranspose_CP_0_elements(378)); -- 
    rr_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(378), ack => type_cast_1224_inst_req_0); -- 
    cr_2840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(378), ack => type_cast_1224_inst_req_1); -- 
    -- CP-element group 379:  transition  place  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	457 
    -- CP-element group 379:  members (5) 
      -- CP-element group 379: 	 branch_block_stmt_25/if_stmt_1197_else_link/$exit
      -- CP-element group 379: 	 branch_block_stmt_25/if_stmt_1197_else_link/else_choice_transition
      -- CP-element group 379: 	 branch_block_stmt_25/forx_xend273_forx_xend428
      -- CP-element group 379: 	 branch_block_stmt_25/forx_xend273_forx_xend428_PhiReq/$entry
      -- CP-element group 379: 	 branch_block_stmt_25/forx_xend273_forx_xend428_PhiReq/$exit
      -- 
    else_choice_transition_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1197_branch_ack_0, ack => convTranspose_CP_0_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: successors 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Sample/ra
      -- 
    ra_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1224_inst_ack_0, ack => convTranspose_CP_0_elements(380)); -- 
    -- CP-element group 381:  transition  place  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	378 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	451 
    -- CP-element group 381:  members (9) 
      -- CP-element group 381: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238__exit__
      -- CP-element group 381: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356
      -- CP-element group 381: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/$entry
      -- CP-element group 381: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/phi_stmt_1241/$entry
      -- CP-element group 381: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/$entry
      -- CP-element group 381: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/$exit
      -- CP-element group 381: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_25/assign_stmt_1209_to_assign_stmt_1238/type_cast_1224_Update/ca
      -- 
    ca_2841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1224_inst_ack_1, ack => convTranspose_CP_0_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	456 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	427 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_sample_complete
      -- CP-element group 382: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Sample/ack
      -- 
    ack_2870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1253_index_offset_ack_0, ack => convTranspose_CP_0_elements(382)); -- 
    -- CP-element group 383:  transition  input  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	456 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (11) 
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_root_address_calculated
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_offset_calculated
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Update/ack
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_base_plus_offset/$entry
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_base_plus_offset/$exit
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_base_plus_offset/sum_rename_req
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_base_plus_offset/sum_rename_ack
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_request/$entry
      -- CP-element group 383: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_request/req
      -- 
    ack_2875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1253_index_offset_ack_1, ack => convTranspose_CP_0_elements(383)); -- 
    req_2884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(383), ack => addr_of_1254_final_reg_req_0); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_request/$exit
      -- CP-element group 384: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_request/ack
      -- 
    ack_2885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1254_final_reg_ack_0, ack => convTranspose_CP_0_elements(384)); -- 
    -- CP-element group 385:  join  fork  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	456 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (24) 
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_complete/$exit
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_complete/ack
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_address_calculated
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_word_address_calculated
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_root_address_calculated
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_address_resized
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_addr_resize/$entry
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_addr_resize/$exit
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_addr_resize/base_resize_req
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_addr_resize/base_resize_ack
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_plus_offset/$entry
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_plus_offset/$exit
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_plus_offset/sum_rename_req
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_base_plus_offset/sum_rename_ack
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_word_addrgen/$entry
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_word_addrgen/$exit
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_word_addrgen/root_register_req
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_word_addrgen/root_register_ack
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/word_access_start/$entry
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/word_access_start/word_0/$entry
      -- CP-element group 385: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/word_access_start/word_0/rr
      -- 
    ack_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1254_final_reg_ack_1, ack => convTranspose_CP_0_elements(385)); -- 
    rr_2923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(385), ack => ptr_deref_1258_load_0_req_0); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (5) 
      -- CP-element group 386: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/word_access_start/$exit
      -- CP-element group 386: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/word_access_start/word_0/$exit
      -- CP-element group 386: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Sample/word_access_start/word_0/ra
      -- 
    ra_2924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1258_load_0_ack_0, ack => convTranspose_CP_0_elements(386)); -- 
    -- CP-element group 387:  fork  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	456 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387: 	390 
    -- CP-element group 387: 	392 
    -- CP-element group 387: 	394 
    -- CP-element group 387: 	396 
    -- CP-element group 387: 	398 
    -- CP-element group 387: 	400 
    -- CP-element group 387: 	402 
    -- CP-element group 387:  members (33) 
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/word_access_complete/$exit
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/word_access_complete/word_0/$exit
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/word_access_complete/word_0/ca
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/ptr_deref_1258_Merge/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/ptr_deref_1258_Merge/$exit
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/ptr_deref_1258_Merge/merge_req
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/ptr_deref_1258_Merge/merge_ack
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_sample_start_
      -- 
    ca_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1258_load_0_ack_1, ack => convTranspose_CP_0_elements(387)); -- 
    rr_2948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1262_inst_req_0); -- 
    rr_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1272_inst_req_0); -- 
    rr_2976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1282_inst_req_0); -- 
    rr_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1292_inst_req_0); -- 
    rr_3004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1302_inst_req_0); -- 
    rr_3018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1312_inst_req_0); -- 
    rr_3032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1322_inst_req_0); -- 
    rr_3046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(387), ack => type_cast_1332_inst_req_0); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Sample/ra
      -- 
    ra_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1262_inst_ack_0, ack => convTranspose_CP_0_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	456 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	424 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Update/ca
      -- 
    ca_2954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1262_inst_ack_1, ack => convTranspose_CP_0_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	387 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Sample/ra
      -- 
    ra_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1272_inst_ack_0, ack => convTranspose_CP_0_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	456 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	421 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Update/ca
      -- 
    ca_2968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1272_inst_ack_1, ack => convTranspose_CP_0_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	387 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Sample/ra
      -- 
    ra_2977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1282_inst_ack_0, ack => convTranspose_CP_0_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	456 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	418 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Update/ca
      -- 
    ca_2982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1282_inst_ack_1, ack => convTranspose_CP_0_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	387 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Sample/ra
      -- 
    ra_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1292_inst_ack_0, ack => convTranspose_CP_0_elements(394)); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	456 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	415 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_update_completed_
      -- CP-element group 395: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Update/ca
      -- 
    ca_2996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1292_inst_ack_1, ack => convTranspose_CP_0_elements(395)); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	387 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_sample_completed_
      -- CP-element group 396: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Sample/ra
      -- 
    ra_3005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_0, ack => convTranspose_CP_0_elements(396)); -- 
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	456 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	412 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_update_completed_
      -- CP-element group 397: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Update/ca
      -- 
    ca_3010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_1, ack => convTranspose_CP_0_elements(397)); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	387 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Sample/ra
      -- CP-element group 398: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_sample_completed_
      -- 
    ra_3019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_0, ack => convTranspose_CP_0_elements(398)); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	456 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	409 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Update/ca
      -- CP-element group 399: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_update_completed_
      -- 
    ca_3024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_1, ack => convTranspose_CP_0_elements(399)); -- 
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	387 
    -- CP-element group 400: successors 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_sample_completed_
      -- CP-element group 400: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Sample/ra
      -- 
    ra_3033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1322_inst_ack_0, ack => convTranspose_CP_0_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	456 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	406 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_update_completed_
      -- CP-element group 401: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Update/ca
      -- CP-element group 401: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Update/$exit
      -- 
    ca_3038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1322_inst_ack_1, ack => convTranspose_CP_0_elements(401)); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	387 
    -- CP-element group 402: successors 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Sample/$exit
      -- CP-element group 402: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Sample/ra
      -- CP-element group 402: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_sample_completed_
      -- 
    ra_3047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_0, ack => convTranspose_CP_0_elements(402)); -- 
    -- CP-element group 403:  transition  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	456 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (6) 
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_update_completed_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Sample/req
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Update/ca
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Update/$exit
      -- 
    ca_3052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_1, ack => convTranspose_CP_0_elements(403)); -- 
    req_3060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(403), ack => WPIPE_ConvTranspose_output_pipe_1334_inst_req_0); -- 
    -- CP-element group 404:  transition  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (6) 
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Update/req
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Sample/ack
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_update_start_
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_sample_completed_
      -- 
    ack_3061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1334_inst_ack_0, ack => convTranspose_CP_0_elements(404)); -- 
    req_3065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(404), ack => WPIPE_ConvTranspose_output_pipe_1334_inst_req_1); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Update/ack
      -- CP-element group 405: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1334_update_completed_
      -- 
    ack_3066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1334_inst_ack_1, ack => convTranspose_CP_0_elements(405)); -- 
    -- CP-element group 406:  join  transition  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	401 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Sample/req
      -- CP-element group 406: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_sample_start_
      -- 
    req_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1337_inst_req_0); -- 
    convTranspose_cp_element_group_406: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_406"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(401) & convTranspose_CP_0_elements(405);
      gj_convTranspose_cp_element_group_406 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(406), clk => clk, reset => reset); --
    end block;
    -- CP-element group 407:  transition  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (6) 
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Update/req
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Sample/ack
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_update_start_
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_sample_completed_
      -- 
    ack_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1337_inst_ack_0, ack => convTranspose_CP_0_elements(407)); -- 
    req_3079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(407), ack => WPIPE_ConvTranspose_output_pipe_1337_inst_req_1); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Update/ack
      -- CP-element group 408: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1337_update_completed_
      -- 
    ack_3080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1337_inst_ack_1, ack => convTranspose_CP_0_elements(408)); -- 
    -- CP-element group 409:  join  transition  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	399 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Sample/req
      -- CP-element group 409: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Sample/$entry
      -- CP-element group 409: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_sample_start_
      -- 
    req_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1340_inst_req_0); -- 
    convTranspose_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(399) & convTranspose_CP_0_elements(408);
      gj_convTranspose_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  transition  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (6) 
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Update/req
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Sample/ack
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_update_start_
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_sample_completed_
      -- 
    ack_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1340_inst_ack_0, ack => convTranspose_CP_0_elements(410)); -- 
    req_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(410), ack => WPIPE_ConvTranspose_output_pipe_1340_inst_req_1); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Update/ack
      -- CP-element group 411: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1340_update_completed_
      -- 
    ack_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1340_inst_ack_1, ack => convTranspose_CP_0_elements(411)); -- 
    -- CP-element group 412:  join  transition  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	397 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Sample/$entry
      -- CP-element group 412: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_sample_start_
      -- CP-element group 412: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Sample/req
      -- 
    req_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1343_inst_req_0); -- 
    convTranspose_cp_element_group_412: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_412"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(397) & convTranspose_CP_0_elements(411);
      gj_convTranspose_cp_element_group_412 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(412), clk => clk, reset => reset); --
    end block;
    -- CP-element group 413:  transition  input  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (6) 
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_sample_completed_
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Sample/ack
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Update/$entry
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Sample/$exit
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_update_start_
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Update/req
      -- 
    ack_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1343_inst_ack_0, ack => convTranspose_CP_0_elements(413)); -- 
    req_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(413), ack => WPIPE_ConvTranspose_output_pipe_1343_inst_req_1); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_update_completed_
      -- CP-element group 414: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Update/$exit
      -- CP-element group 414: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1343_Update/ack
      -- 
    ack_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1343_inst_ack_1, ack => convTranspose_CP_0_elements(414)); -- 
    -- CP-element group 415:  join  transition  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	395 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_sample_start_
      -- CP-element group 415: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Sample/req
      -- 
    req_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1346_inst_req_0); -- 
    convTranspose_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(395) & convTranspose_CP_0_elements(414);
      gj_convTranspose_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  transition  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (6) 
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_sample_completed_
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_update_start_
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Update/req
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Update/$entry
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Sample/$exit
      -- 
    ack_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1346_inst_ack_0, ack => convTranspose_CP_0_elements(416)); -- 
    req_3121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(416), ack => WPIPE_ConvTranspose_output_pipe_1346_inst_req_1); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1346_Update/$exit
      -- 
    ack_3122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1346_inst_ack_1, ack => convTranspose_CP_0_elements(417)); -- 
    -- CP-element group 418:  join  transition  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	393 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_sample_start_
      -- 
    req_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(418), ack => WPIPE_ConvTranspose_output_pipe_1349_inst_req_0); -- 
    convTranspose_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(393) & convTranspose_CP_0_elements(417);
      gj_convTranspose_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  transition  input  output  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (6) 
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Update/req
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Update/$entry
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Sample/ack
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_update_start_
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_sample_completed_
      -- 
    ack_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1349_inst_ack_0, ack => convTranspose_CP_0_elements(419)); -- 
    req_3135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(419), ack => WPIPE_ConvTranspose_output_pipe_1349_inst_req_1); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Update/ack
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1349_update_completed_
      -- 
    ack_3136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1349_inst_ack_1, ack => convTranspose_CP_0_elements(420)); -- 
    -- CP-element group 421:  join  transition  output  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	391 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Sample/req
      -- CP-element group 421: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Sample/$entry
      -- CP-element group 421: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_sample_start_
      -- 
    req_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(421), ack => WPIPE_ConvTranspose_output_pipe_1352_inst_req_0); -- 
    convTranspose_cp_element_group_421: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_421"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(391) & convTranspose_CP_0_elements(420);
      gj_convTranspose_cp_element_group_421 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(421), clk => clk, reset => reset); --
    end block;
    -- CP-element group 422:  transition  input  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (6) 
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Update/req
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Update/$entry
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Sample/ack
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Sample/$exit
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_update_start_
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_sample_completed_
      -- 
    ack_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1352_inst_ack_0, ack => convTranspose_CP_0_elements(422)); -- 
    req_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(422), ack => WPIPE_ConvTranspose_output_pipe_1352_inst_req_1); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Update/ack
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_Update/$exit
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1352_update_completed_
      -- 
    ack_3150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1352_inst_ack_1, ack => convTranspose_CP_0_elements(423)); -- 
    -- CP-element group 424:  join  transition  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	389 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Sample/req
      -- CP-element group 424: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_sample_start_
      -- 
    req_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(424), ack => WPIPE_ConvTranspose_output_pipe_1355_inst_req_0); -- 
    convTranspose_cp_element_group_424: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_424"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(389) & convTranspose_CP_0_elements(423);
      gj_convTranspose_cp_element_group_424 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(424), clk => clk, reset => reset); --
    end block;
    -- CP-element group 425:  transition  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (6) 
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Update/req
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Update/$entry
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Sample/ack
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_update_start_
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_sample_completed_
      -- 
    ack_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1355_inst_ack_0, ack => convTranspose_CP_0_elements(425)); -- 
    req_3163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(425), ack => WPIPE_ConvTranspose_output_pipe_1355_inst_req_1); -- 
    -- CP-element group 426:  transition  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Update/ack
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/WPIPE_ConvTranspose_output_pipe_1355_update_completed_
      -- 
    ack_3164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1355_inst_ack_1, ack => convTranspose_CP_0_elements(426)); -- 
    -- CP-element group 427:  branch  join  transition  place  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	382 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427: 	429 
    -- CP-element group 427:  members (10) 
      -- CP-element group 427: 	 branch_block_stmt_25/if_stmt_1369_eval_test/$exit
      -- CP-element group 427: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368__exit__
      -- CP-element group 427: 	 branch_block_stmt_25/if_stmt_1369__entry__
      -- CP-element group 427: 	 branch_block_stmt_25/if_stmt_1369_if_link/$entry
      -- CP-element group 427: 	 branch_block_stmt_25/if_stmt_1369_eval_test/branch_req
      -- CP-element group 427: 	 branch_block_stmt_25/if_stmt_1369_eval_test/$entry
      -- CP-element group 427: 	 branch_block_stmt_25/if_stmt_1369_else_link/$entry
      -- CP-element group 427: 	 branch_block_stmt_25/if_stmt_1369_dead_link/$entry
      -- CP-element group 427: 	 branch_block_stmt_25/R_exitcond1_1370_place
      -- CP-element group 427: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/$exit
      -- 
    branch_req_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(427), ack => if_stmt_1369_branch_req_0); -- 
    convTranspose_cp_element_group_427: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_427"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(382) & convTranspose_CP_0_elements(426);
      gj_convTranspose_cp_element_group_427 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(427), clk => clk, reset => reset); --
    end block;
    -- CP-element group 428:  merge  transition  place  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	457 
    -- CP-element group 428:  members (13) 
      -- CP-element group 428: 	 branch_block_stmt_25/merge_stmt_1375__exit__
      -- CP-element group 428: 	 branch_block_stmt_25/forx_xend428x_xloopexit_forx_xend428
      -- CP-element group 428: 	 branch_block_stmt_25/if_stmt_1369_if_link/if_choice_transition
      -- CP-element group 428: 	 branch_block_stmt_25/if_stmt_1369_if_link/$exit
      -- CP-element group 428: 	 branch_block_stmt_25/forx_xbody356_forx_xend428x_xloopexit
      -- CP-element group 428: 	 branch_block_stmt_25/forx_xbody356_forx_xend428x_xloopexit_PhiReq/$entry
      -- CP-element group 428: 	 branch_block_stmt_25/forx_xbody356_forx_xend428x_xloopexit_PhiReq/$exit
      -- CP-element group 428: 	 branch_block_stmt_25/merge_stmt_1375_PhiReqMerge
      -- CP-element group 428: 	 branch_block_stmt_25/merge_stmt_1375_PhiAck/$entry
      -- CP-element group 428: 	 branch_block_stmt_25/merge_stmt_1375_PhiAck/$exit
      -- CP-element group 428: 	 branch_block_stmt_25/merge_stmt_1375_PhiAck/dummy
      -- CP-element group 428: 	 branch_block_stmt_25/forx_xend428x_xloopexit_forx_xend428_PhiReq/$entry
      -- CP-element group 428: 	 branch_block_stmt_25/forx_xend428x_xloopexit_forx_xend428_PhiReq/$exit
      -- 
    if_choice_transition_3177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1369_branch_ack_1, ack => convTranspose_CP_0_elements(428)); -- 
    -- CP-element group 429:  fork  transition  place  input  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	452 
    -- CP-element group 429: 	453 
    -- CP-element group 429:  members (12) 
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356
      -- CP-element group 429: 	 branch_block_stmt_25/if_stmt_1369_else_link/else_choice_transition
      -- CP-element group 429: 	 branch_block_stmt_25/if_stmt_1369_else_link/$exit
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Update/cr
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Update/$entry
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/$entry
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/$entry
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/$entry
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/$entry
      -- CP-element group 429: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/$entry
      -- 
    else_choice_transition_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1369_branch_ack_0, ack => convTranspose_CP_0_elements(429)); -- 
    cr_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(429), ack => type_cast_1247_inst_req_1); -- 
    rr_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(429), ack => type_cast_1247_inst_req_0); -- 
    -- CP-element group 430:  merge  branch  transition  place  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	120 
    -- CP-element group 430: 	165 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	121 
    -- CP-element group 430: 	122 
    -- CP-element group 430:  members (17) 
      -- CP-element group 430: 	 branch_block_stmt_25/merge_stmt_417__exit__
      -- CP-element group 430: 	 branch_block_stmt_25/assign_stmt_423__entry__
      -- CP-element group 430: 	 branch_block_stmt_25/assign_stmt_423__exit__
      -- CP-element group 430: 	 branch_block_stmt_25/if_stmt_424__entry__
      -- CP-element group 430: 	 branch_block_stmt_25/merge_stmt_417_PhiReqMerge
      -- CP-element group 430: 	 branch_block_stmt_25/assign_stmt_423/$entry
      -- CP-element group 430: 	 branch_block_stmt_25/assign_stmt_423/$exit
      -- CP-element group 430: 	 branch_block_stmt_25/if_stmt_424_dead_link/$entry
      -- CP-element group 430: 	 branch_block_stmt_25/if_stmt_424_eval_test/$entry
      -- CP-element group 430: 	 branch_block_stmt_25/if_stmt_424_eval_test/$exit
      -- CP-element group 430: 	 branch_block_stmt_25/if_stmt_424_eval_test/branch_req
      -- CP-element group 430: 	 branch_block_stmt_25/R_cmp194437_425_place
      -- CP-element group 430: 	 branch_block_stmt_25/if_stmt_424_if_link/$entry
      -- CP-element group 430: 	 branch_block_stmt_25/if_stmt_424_else_link/$entry
      -- CP-element group 430: 	 branch_block_stmt_25/merge_stmt_417_PhiAck/$entry
      -- CP-element group 430: 	 branch_block_stmt_25/merge_stmt_417_PhiAck/$exit
      -- CP-element group 430: 	 branch_block_stmt_25/merge_stmt_417_PhiAck/dummy
      -- 
    branch_req_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(430), ack => if_stmt_424_branch_req_0); -- 
    convTranspose_CP_0_elements(430) <= OrReduce(convTranspose_CP_0_elements(120) & convTranspose_CP_0_elements(165));
    -- CP-element group 431:  transition  output  delay-element  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	124 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	435 
    -- CP-element group 431:  members (5) 
      -- CP-element group 431: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_req
      -- CP-element group 431: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_466_konst_delay_trans
      -- CP-element group 431: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/$exit
      -- CP-element group 431: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/phi_stmt_462/$exit
      -- CP-element group 431: 	 branch_block_stmt_25/bbx_xnph443_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_462_req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_462_req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(431), ack => phi_stmt_462_req_0); -- 
    -- Element group convTranspose_CP_0_elements(431) is a control-delay.
    cp_element_431_delay: control_delay_element  generic map(name => " 431_delay", delay_value => 1)  port map(req => convTranspose_CP_0_elements(124), ack => convTranspose_CP_0_elements(431), clk => clk, reset =>reset);
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	166 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	434 
    -- CP-element group 432:  members (2) 
      -- CP-element group 432: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Sample/ra
      -- CP-element group 432: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Sample/$exit
      -- 
    ra_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_468_inst_ack_0, ack => convTranspose_CP_0_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	166 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (2) 
      -- CP-element group 433: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Update/ca
      -- CP-element group 433: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/Update/$exit
      -- 
    ca_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_468_inst_ack_1, ack => convTranspose_CP_0_elements(433)); -- 
    -- CP-element group 434:  join  transition  output  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	432 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (6) 
      -- CP-element group 434: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_req
      -- CP-element group 434: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/SplitProtocol/$exit
      -- CP-element group 434: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/type_cast_468/$exit
      -- CP-element group 434: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/phi_stmt_462_sources/$exit
      -- CP-element group 434: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_462/$exit
      -- CP-element group 434: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_462_req_3255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_462_req_3255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(434), ack => phi_stmt_462_req_1); -- 
    convTranspose_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(432) & convTranspose_CP_0_elements(433);
      gj_convTranspose_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  merge  transition  place  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	431 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (2) 
      -- CP-element group 435: 	 branch_block_stmt_25/merge_stmt_461_PhiReqMerge
      -- CP-element group 435: 	 branch_block_stmt_25/merge_stmt_461_PhiAck/$entry
      -- 
    convTranspose_CP_0_elements(435) <= OrReduce(convTranspose_CP_0_elements(431) & convTranspose_CP_0_elements(434));
    -- CP-element group 436:  fork  transition  place  input  output  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	125 
    -- CP-element group 436: 	126 
    -- CP-element group 436: 	128 
    -- CP-element group 436: 	129 
    -- CP-element group 436: 	132 
    -- CP-element group 436: 	136 
    -- CP-element group 436: 	140 
    -- CP-element group 436: 	144 
    -- CP-element group 436: 	148 
    -- CP-element group 436: 	152 
    -- CP-element group 436: 	156 
    -- CP-element group 436: 	160 
    -- CP-element group 436: 	163 
    -- CP-element group 436:  members (56) 
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_sample_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_complete/req
      -- CP-element group 436: 	 branch_block_stmt_25/merge_stmt_461__exit__
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624__entry__
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Sample/rr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_513_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/RPIPE_ConvTranspose_input_pipe_478_Sample/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/word_access_complete/word_0/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_585_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/word_access_complete/word_0/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/word_access_complete/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/ptr_deref_611_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_495_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_531_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_603_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_549_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_482_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_complete/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/type_cast_567_Update/cr
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/addr_of_475_update_start_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_resized_1
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_scaled_1
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_computed_1
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_resize_1/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_resize_1/$exit
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_resize_1/index_resize_req
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_resize_1/index_resize_ack
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_scale_1/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_scale_1/$exit
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_scale_1/scale_rename_req
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_index_scale_1/scale_rename_ack
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_update_start
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Sample/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Sample/req
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_476_to_assign_stmt_624/array_obj_ref_474_final_index_sum_regn_Update/req
      -- CP-element group 436: 	 branch_block_stmt_25/merge_stmt_461_PhiAck/phi_stmt_462_ack
      -- CP-element group 436: 	 branch_block_stmt_25/merge_stmt_461_PhiAck/$exit
      -- 
    phi_stmt_462_ack_3260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_462_ack_0, ack => convTranspose_CP_0_elements(436)); -- 
    req_964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => addr_of_475_final_reg_req_1); -- 
    cr_1048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_513_inst_req_1); -- 
    rr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => RPIPE_ConvTranspose_input_pipe_478_inst_req_0); -- 
    cr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_531_inst_req_1); -- 
    cr_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_585_inst_req_1); -- 
    cr_1020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_495_inst_req_1); -- 
    cr_1188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_603_inst_req_1); -- 
    cr_992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_482_inst_req_1); -- 
    cr_1238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => ptr_deref_611_store_0_req_1); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_549_inst_req_1); -- 
    cr_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => type_cast_567_inst_req_1); -- 
    req_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => array_obj_ref_474_index_offset_req_0); -- 
    req_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(436), ack => array_obj_ref_474_index_offset_req_1); -- 
    -- CP-element group 437:  transition  output  delay-element  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	168 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	441 
    -- CP-element group 437:  members (5) 
      -- CP-element group 437: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_675_konst_delay_trans
      -- CP-element group 437: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_req
      -- CP-element group 437: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/$exit
      -- CP-element group 437: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/phi_stmt_669/$exit
      -- CP-element group 437: 	 branch_block_stmt_25/bbx_xnph439_forx_xbody196_PhiReq/$exit
      -- 
    phi_stmt_669_req_3283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_669_req_3283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(437), ack => phi_stmt_669_req_1); -- 
    -- Element group convTranspose_CP_0_elements(437) is a control-delay.
    cp_element_437_delay: control_delay_element  generic map(name => " 437_delay", delay_value => 1)  port map(req => convTranspose_CP_0_elements(168), ack => convTranspose_CP_0_elements(437), clk => clk, reset =>reset);
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	210 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	440 
    -- CP-element group 438:  members (2) 
      -- CP-element group 438: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Sample/ra
      -- CP-element group 438: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Sample/$exit
      -- 
    ra_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_672_inst_ack_0, ack => convTranspose_CP_0_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	210 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (2) 
      -- CP-element group 439: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Update/ca
      -- CP-element group 439: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/Update/$exit
      -- 
    ca_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_672_inst_ack_1, ack => convTranspose_CP_0_elements(439)); -- 
    -- CP-element group 440:  join  transition  output  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	441 
    -- CP-element group 440:  members (6) 
      -- CP-element group 440: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/$exit
      -- CP-element group 440: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/$exit
      -- CP-element group 440: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 440: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/$exit
      -- CP-element group 440: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_sources/type_cast_672/SplitProtocol/$exit
      -- CP-element group 440: 	 branch_block_stmt_25/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_669/phi_stmt_669_req
      -- 
    phi_stmt_669_req_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_669_req_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(440), ack => phi_stmt_669_req_0); -- 
    convTranspose_cp_element_group_440: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_440"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(438) & convTranspose_CP_0_elements(439);
      gj_convTranspose_cp_element_group_440 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(440), clk => clk, reset => reset); --
    end block;
    -- CP-element group 441:  merge  transition  place  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	437 
    -- CP-element group 441: 	440 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441:  members (2) 
      -- CP-element group 441: 	 branch_block_stmt_25/merge_stmt_668_PhiReqMerge
      -- CP-element group 441: 	 branch_block_stmt_25/merge_stmt_668_PhiAck/$entry
      -- 
    convTranspose_CP_0_elements(441) <= OrReduce(convTranspose_CP_0_elements(437) & convTranspose_CP_0_elements(440));
    -- CP-element group 442:  fork  transition  place  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	169 
    -- CP-element group 442: 	170 
    -- CP-element group 442: 	172 
    -- CP-element group 442: 	173 
    -- CP-element group 442: 	176 
    -- CP-element group 442: 	180 
    -- CP-element group 442: 	184 
    -- CP-element group 442: 	188 
    -- CP-element group 442: 	192 
    -- CP-element group 442: 	196 
    -- CP-element group 442: 	200 
    -- CP-element group 442: 	204 
    -- CP-element group 442: 	207 
    -- CP-element group 442:  members (56) 
      -- CP-element group 442: 	 branch_block_stmt_25/merge_stmt_668__exit__
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831__entry__
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_resize_1/$exit
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Sample/rr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_resize_1/index_resize_ack
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_resize_1/index_resize_req
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/RPIPE_ConvTranspose_input_pipe_685_sample_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_resize_1/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_computed_1
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_scaled_1
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_resized_1
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_complete/req
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/addr_of_682_complete/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_720_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/merge_stmt_668_PhiAck/phi_stmt_669_ack
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Update/req
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Sample/req
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_702_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_final_index_sum_regn_update_start
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_689_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_scale_1/scale_rename_ack
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_scale_1/scale_rename_req
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_scale_1/$exit
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/array_obj_ref_681_index_scale_1/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_738_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_756_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_774_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/merge_stmt_668_PhiAck/$exit
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_792_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/type_cast_810_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_update_start_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/word_access_complete/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/word_access_complete/word_0/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_683_to_assign_stmt_831/ptr_deref_818_Update/word_access_complete/word_0/cr
      -- 
    phi_stmt_669_ack_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_669_ack_0, ack => convTranspose_CP_0_elements(442)); -- 
    rr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => RPIPE_ConvTranspose_input_pipe_685_inst_req_0); -- 
    cr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_702_inst_req_1); -- 
    req_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => addr_of_682_final_reg_req_1); -- 
    cr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_720_inst_req_1); -- 
    req_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => array_obj_ref_681_index_offset_req_1); -- 
    req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => array_obj_ref_681_index_offset_req_0); -- 
    cr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_689_inst_req_1); -- 
    cr_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_738_inst_req_1); -- 
    cr_1463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_756_inst_req_1); -- 
    cr_1491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_774_inst_req_1); -- 
    cr_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_792_inst_req_1); -- 
    cr_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => type_cast_810_inst_req_1); -- 
    cr_1597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(442), ack => ptr_deref_818_store_0_req_1); -- 
    -- CP-element group 443:  merge  fork  transition  place  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	122 
    -- CP-element group 443: 	209 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	211 
    -- CP-element group 443: 	212 
    -- CP-element group 443: 	213 
    -- CP-element group 443: 	214 
    -- CP-element group 443: 	215 
    -- CP-element group 443: 	216 
    -- CP-element group 443:  members (25) 
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_840__exit__
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868__entry__
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_840_PhiReqMerge
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_update_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Sample/rr
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_843_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_update_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Sample/rr
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_847_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_update_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Sample/rr
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_844_to_assign_stmt_868/type_cast_851_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_840_PhiAck/dummy
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_840_PhiAck/$exit
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_840_PhiAck/$entry
      -- 
    rr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(443), ack => type_cast_843_inst_req_0); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(443), ack => type_cast_843_inst_req_1); -- 
    rr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(443), ack => type_cast_847_inst_req_0); -- 
    cr_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(443), ack => type_cast_847_inst_req_1); -- 
    rr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(443), ack => type_cast_851_inst_req_0); -- 
    cr_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(443), ack => type_cast_851_inst_req_1); -- 
    convTranspose_CP_0_elements(443) <= OrReduce(convTranspose_CP_0_elements(122) & convTranspose_CP_0_elements(209));
    -- CP-element group 444:  transition  output  delay-element  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	221 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	448 
    -- CP-element group 444:  members (5) 
      -- CP-element group 444: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/$exit
      -- CP-element group 444: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919_konst_delay_trans
      -- CP-element group 444: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_req
      -- CP-element group 444: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/phi_stmt_913/$exit
      -- CP-element group 444: 	 branch_block_stmt_25/bbx_xnph435_forx_xbody266_PhiReq/$exit
      -- 
    phi_stmt_913_req_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_913_req_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(444), ack => phi_stmt_913_req_1); -- 
    -- Element group convTranspose_CP_0_elements(444) is a control-delay.
    cp_element_444_delay: control_delay_element  generic map(name => " 444_delay", delay_value => 1)  port map(req => convTranspose_CP_0_elements(221), ack => convTranspose_CP_0_elements(444), clk => clk, reset =>reset);
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	230 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	447 
    -- CP-element group 445:  members (2) 
      -- CP-element group 445: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Sample/$exit
      -- CP-element group 445: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Sample/ra
      -- 
    ra_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_0, ack => convTranspose_CP_0_elements(445)); -- 
    -- CP-element group 446:  transition  input  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	230 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (2) 
      -- CP-element group 446: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Update/ca
      -- CP-element group 446: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/Update/$exit
      -- 
    ca_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_1, ack => convTranspose_CP_0_elements(446)); -- 
    -- CP-element group 447:  join  transition  output  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	445 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (6) 
      -- CP-element group 447: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/$exit
      -- CP-element group 447: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 447: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/SplitProtocol/$exit
      -- CP-element group 447: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_916/$exit
      -- CP-element group 447: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/phi_stmt_913_req
      -- CP-element group 447: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_913/$exit
      -- 
    phi_stmt_913_req_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_913_req_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(447), ack => phi_stmt_913_req_0); -- 
    convTranspose_cp_element_group_447: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_447"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(445) & convTranspose_CP_0_elements(446);
      gj_convTranspose_cp_element_group_447 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(447), clk => clk, reset => reset); --
    end block;
    -- CP-element group 448:  merge  transition  place  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	444 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (2) 
      -- CP-element group 448: 	 branch_block_stmt_25/merge_stmt_912_PhiReqMerge
      -- CP-element group 448: 	 branch_block_stmt_25/merge_stmt_912_PhiAck/$entry
      -- 
    convTranspose_CP_0_elements(448) <= OrReduce(convTranspose_CP_0_elements(444) & convTranspose_CP_0_elements(447));
    -- CP-element group 449:  fork  transition  place  input  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	222 
    -- CP-element group 449: 	223 
    -- CP-element group 449: 	225 
    -- CP-element group 449: 	227 
    -- CP-element group 449:  members (29) 
      -- CP-element group 449: 	 branch_block_stmt_25/merge_stmt_912__exit__
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943__entry__
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_update_start_
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_resized_1
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_scaled_1
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_computed_1
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_resize_1/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_resize_1/$exit
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_resize_1/index_resize_req
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_resize_1/index_resize_ack
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_scale_1/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_scale_1/$exit
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_scale_1/scale_rename_req
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_index_scale_1/scale_rename_ack
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_update_start
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Sample/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Sample/req
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/array_obj_ref_925_final_index_sum_regn_Update/req
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_complete/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/addr_of_926_complete/req
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_update_start_
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/word_access_complete/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/word_access_complete/word_0/$entry
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_927_to_assign_stmt_943/ptr_deref_929_Update/word_access_complete/word_0/cr
      -- CP-element group 449: 	 branch_block_stmt_25/merge_stmt_912_PhiAck/phi_stmt_913_ack
      -- CP-element group 449: 	 branch_block_stmt_25/merge_stmt_912_PhiAck/$exit
      -- 
    phi_stmt_913_ack_3391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_913_ack_0, ack => convTranspose_CP_0_elements(449)); -- 
    req_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(449), ack => array_obj_ref_925_index_offset_req_0); -- 
    req_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(449), ack => array_obj_ref_925_index_offset_req_1); -- 
    req_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(449), ack => addr_of_926_final_reg_req_1); -- 
    cr_1796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(449), ack => ptr_deref_929_store_0_req_1); -- 
    -- CP-element group 450:  merge  transition  place  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	219 
    -- CP-element group 450: 	229 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	231 
    -- CP-element group 450:  members (10) 
      -- CP-element group 450: 	 branch_block_stmt_25/merge_stmt_952__exit__
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961__entry__
      -- CP-element group 450: 	 branch_block_stmt_25/merge_stmt_952_PhiReqMerge
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_sample_start_
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Sample/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_957_to_assign_stmt_961/WPIPE_ConvTranspose_output_pipe_954_Sample/req
      -- CP-element group 450: 	 branch_block_stmt_25/merge_stmt_952_PhiAck/dummy
      -- CP-element group 450: 	 branch_block_stmt_25/merge_stmt_952_PhiAck/$exit
      -- CP-element group 450: 	 branch_block_stmt_25/merge_stmt_952_PhiAck/$entry
      -- 
    req_1827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(450), ack => WPIPE_ConvTranspose_output_pipe_954_inst_req_0); -- 
    convTranspose_CP_0_elements(450) <= OrReduce(convTranspose_CP_0_elements(219) & convTranspose_CP_0_elements(229));
    -- CP-element group 451:  transition  output  delay-element  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	381 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	455 
    -- CP-element group 451:  members (5) 
      -- CP-element group 451: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_req
      -- CP-element group 451: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1245_konst_delay_trans
      -- CP-element group 451: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/$exit
      -- CP-element group 451: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/phi_stmt_1241/$exit
      -- CP-element group 451: 	 branch_block_stmt_25/bbx_xnph_forx_xbody356_PhiReq/$exit
      -- 
    phi_stmt_1241_req_3437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1241_req_3437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(451), ack => phi_stmt_1241_req_0); -- 
    -- Element group convTranspose_CP_0_elements(451) is a control-delay.
    cp_element_451_delay: control_delay_element  generic map(name => " 451_delay", delay_value => 1)  port map(req => convTranspose_CP_0_elements(381), ack => convTranspose_CP_0_elements(451), clk => clk, reset =>reset);
    -- CP-element group 452:  transition  input  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	429 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	454 
    -- CP-element group 452:  members (2) 
      -- CP-element group 452: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Sample/ra
      -- CP-element group 452: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Sample/$exit
      -- 
    ra_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_0, ack => convTranspose_CP_0_elements(452)); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	429 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (2) 
      -- CP-element group 453: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Update/ca
      -- CP-element group 453: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/Update/$exit
      -- 
    ca_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_1, ack => convTranspose_CP_0_elements(453)); -- 
    -- CP-element group 454:  join  transition  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	452 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (6) 
      -- CP-element group 454: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_req
      -- CP-element group 454: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/SplitProtocol/$exit
      -- CP-element group 454: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/type_cast_1247/$exit
      -- CP-element group 454: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/phi_stmt_1241_sources/$exit
      -- CP-element group 454: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/phi_stmt_1241/$exit
      -- CP-element group 454: 	 branch_block_stmt_25/forx_xbody356_forx_xbody356_PhiReq/$exit
      -- 
    phi_stmt_1241_req_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1241_req_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(454), ack => phi_stmt_1241_req_1); -- 
    convTranspose_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_0_elements(452) & convTranspose_CP_0_elements(453);
      gj_convTranspose_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_0_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  merge  transition  place  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	451 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (2) 
      -- CP-element group 455: 	 branch_block_stmt_25/merge_stmt_1240_PhiAck/$entry
      -- CP-element group 455: 	 branch_block_stmt_25/merge_stmt_1240_PhiReqMerge
      -- 
    convTranspose_CP_0_elements(455) <= OrReduce(convTranspose_CP_0_elements(451) & convTranspose_CP_0_elements(454));
    -- CP-element group 456:  fork  transition  place  input  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	382 
    -- CP-element group 456: 	383 
    -- CP-element group 456: 	385 
    -- CP-element group 456: 	387 
    -- CP-element group 456: 	389 
    -- CP-element group 456: 	391 
    -- CP-element group 456: 	393 
    -- CP-element group 456: 	395 
    -- CP-element group 456: 	397 
    -- CP-element group 456: 	399 
    -- CP-element group 456: 	401 
    -- CP-element group 456: 	403 
    -- CP-element group 456:  members (53) 
      -- CP-element group 456: 	 branch_block_stmt_25/merge_stmt_1240__exit__
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368__entry__
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/merge_stmt_1240_PhiAck/phi_stmt_1241_ack
      -- CP-element group 456: 	 branch_block_stmt_25/merge_stmt_1240_PhiAck/$exit
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1322_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1332_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_resized_1
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_scaled_1
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_computed_1
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_resize_1/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_resize_1/$exit
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_resize_1/index_resize_req
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_resize_1/index_resize_ack
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_scale_1/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_scale_1/$exit
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_scale_1/scale_rename_req
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_index_scale_1/scale_rename_ack
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_update_start
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Sample/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Sample/req
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/array_obj_ref_1253_final_index_sum_regn_Update/req
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_complete/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/addr_of_1254_complete/req
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/word_access_complete/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/word_access_complete/word_0/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/ptr_deref_1258_Update/word_access_complete/word_0/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1262_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1272_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1282_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1292_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_update_start_
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1302_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1255_to_assign_stmt_1368/type_cast_1312_update_start_
      -- 
    phi_stmt_1241_ack_3468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1241_ack_0, ack => convTranspose_CP_0_elements(456)); -- 
    cr_3023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1312_inst_req_1); -- 
    cr_3037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1322_inst_req_1); -- 
    cr_3051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1332_inst_req_1); -- 
    req_2869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => array_obj_ref_1253_index_offset_req_0); -- 
    req_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => array_obj_ref_1253_index_offset_req_1); -- 
    req_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => addr_of_1254_final_reg_req_1); -- 
    cr_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => ptr_deref_1258_load_0_req_1); -- 
    cr_2953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1262_inst_req_1); -- 
    cr_2967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1272_inst_req_1); -- 
    cr_2981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1282_inst_req_1); -- 
    cr_2995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1292_inst_req_1); -- 
    cr_3009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_0_elements(456), ack => type_cast_1302_inst_req_1); -- 
    -- CP-element group 457:  merge  transition  place  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	379 
    -- CP-element group 457: 	428 
    -- CP-element group 457: successors 
    -- CP-element group 457:  members (16) 
      -- CP-element group 457: 	 branch_block_stmt_25/branch_block_stmt_25__exit__
      -- CP-element group 457: 	 $exit
      -- CP-element group 457: 	 branch_block_stmt_25/$exit
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1377__exit__
      -- CP-element group 457: 	 branch_block_stmt_25/return__
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1379__exit__
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1377_PhiReqMerge
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1377_PhiAck/$entry
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1377_PhiAck/$exit
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1377_PhiAck/dummy
      -- CP-element group 457: 	 branch_block_stmt_25/return___PhiReq/$entry
      -- CP-element group 457: 	 branch_block_stmt_25/return___PhiReq/$exit
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1379_PhiReqMerge
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1379_PhiAck/$entry
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1379_PhiAck/$exit
      -- CP-element group 457: 	 branch_block_stmt_25/merge_stmt_1379_PhiAck/dummy
      -- 
    convTranspose_CP_0_elements(457) <= OrReduce(convTranspose_CP_0_elements(379) & convTranspose_CP_0_elements(428));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar453_924_resized : std_logic_vector(13 downto 0);
    signal R_indvar453_924_scaled : std_logic_vector(13 downto 0);
    signal R_indvar467_680_resized : std_logic_vector(10 downto 0);
    signal R_indvar467_680_scaled : std_logic_vector(10 downto 0);
    signal R_indvar483_473_resized : std_logic_vector(13 downto 0);
    signal R_indvar483_473_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1252_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1252_scaled : std_logic_vector(13 downto 0);
    signal add108_326 : std_logic_vector(15 downto 0);
    signal add117_351 : std_logic_vector(15 downto 0);
    signal add126_376 : std_logic_vector(15 downto 0);
    signal add12_75 : std_logic_vector(15 downto 0);
    signal add135_401 : std_logic_vector(15 downto 0);
    signal add150_501 : std_logic_vector(63 downto 0);
    signal add156_519 : std_logic_vector(63 downto 0);
    signal add162_537 : std_logic_vector(63 downto 0);
    signal add168_555 : std_logic_vector(63 downto 0);
    signal add174_573 : std_logic_vector(63 downto 0);
    signal add180_591 : std_logic_vector(63 downto 0);
    signal add186_609 : std_logic_vector(63 downto 0);
    signal add206_708 : std_logic_vector(63 downto 0);
    signal add212_726 : std_logic_vector(63 downto 0);
    signal add218_744 : std_logic_vector(63 downto 0);
    signal add21_100 : std_logic_vector(15 downto 0);
    signal add224_762 : std_logic_vector(63 downto 0);
    signal add230_780 : std_logic_vector(63 downto 0);
    signal add236_798 : std_logic_vector(63 downto 0);
    signal add242_816 : std_logic_vector(63 downto 0);
    signal add30_125 : std_logic_vector(15 downto 0);
    signal add39_150 : std_logic_vector(15 downto 0);
    signal add48_175 : std_logic_vector(15 downto 0);
    signal add57_200 : std_logic_vector(15 downto 0);
    signal add74_240 : std_logic_vector(31 downto 0);
    signal add79_245 : std_logic_vector(31 downto 0);
    signal add99_301 : std_logic_vector(15 downto 0);
    signal add_50 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1253_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1253_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1253_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1253_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1253_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1253_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_474_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_474_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_474_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_474_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_474_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_474_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_681_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_681_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_681_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_681_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_681_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_681_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_925_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_925_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_925_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_925_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_925_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_925_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_683 : std_logic_vector(31 downto 0);
    signal arrayidx269_927 : std_logic_vector(31 downto 0);
    signal arrayidx361_1255 : std_logic_vector(31 downto 0);
    signal arrayidx_476 : std_logic_vector(31 downto 0);
    signal call101_304 : std_logic_vector(7 downto 0);
    signal call106_317 : std_logic_vector(7 downto 0);
    signal call10_66 : std_logic_vector(7 downto 0);
    signal call110_329 : std_logic_vector(7 downto 0);
    signal call115_342 : std_logic_vector(7 downto 0);
    signal call119_354 : std_logic_vector(7 downto 0);
    signal call124_367 : std_logic_vector(7 downto 0);
    signal call128_379 : std_logic_vector(7 downto 0);
    signal call133_392 : std_logic_vector(7 downto 0);
    signal call143_479 : std_logic_vector(7 downto 0);
    signal call147_492 : std_logic_vector(7 downto 0);
    signal call14_78 : std_logic_vector(7 downto 0);
    signal call153_510 : std_logic_vector(7 downto 0);
    signal call159_528 : std_logic_vector(7 downto 0);
    signal call165_546 : std_logic_vector(7 downto 0);
    signal call171_564 : std_logic_vector(7 downto 0);
    signal call177_582 : std_logic_vector(7 downto 0);
    signal call183_600 : std_logic_vector(7 downto 0);
    signal call199_686 : std_logic_vector(7 downto 0);
    signal call19_91 : std_logic_vector(7 downto 0);
    signal call203_699 : std_logic_vector(7 downto 0);
    signal call209_717 : std_logic_vector(7 downto 0);
    signal call215_735 : std_logic_vector(7 downto 0);
    signal call221_753 : std_logic_vector(7 downto 0);
    signal call227_771 : std_logic_vector(7 downto 0);
    signal call233_789 : std_logic_vector(7 downto 0);
    signal call239_807 : std_logic_vector(7 downto 0);
    signal call23_103 : std_logic_vector(7 downto 0);
    signal call28_116 : std_logic_vector(7 downto 0);
    signal call2_41 : std_logic_vector(7 downto 0);
    signal call32_128 : std_logic_vector(7 downto 0);
    signal call343_1177 : std_logic_vector(15 downto 0);
    signal call345_1180 : std_logic_vector(15 downto 0);
    signal call347_1183 : std_logic_vector(15 downto 0);
    signal call349_1186 : std_logic_vector(15 downto 0);
    signal call37_141 : std_logic_vector(7 downto 0);
    signal call41_153 : std_logic_vector(7 downto 0);
    signal call46_166 : std_logic_vector(7 downto 0);
    signal call50_178 : std_logic_vector(7 downto 0);
    signal call55_191 : std_logic_vector(7 downto 0);
    signal call5_53 : std_logic_vector(7 downto 0);
    signal call92_279 : std_logic_vector(7 downto 0);
    signal call97_292 : std_logic_vector(7 downto 0);
    signal call_28 : std_logic_vector(7 downto 0);
    signal cmp194437_423 : std_logic_vector(0 downto 0);
    signal cmp264433_868 : std_logic_vector(0 downto 0);
    signal cmp441_408 : std_logic_vector(0 downto 0);
    signal conv104_308 : std_logic_vector(15 downto 0);
    signal conv107_321 : std_logic_vector(15 downto 0);
    signal conv113_333 : std_logic_vector(15 downto 0);
    signal conv116_346 : std_logic_vector(15 downto 0);
    signal conv11_70 : std_logic_vector(15 downto 0);
    signal conv122_358 : std_logic_vector(15 downto 0);
    signal conv125_371 : std_logic_vector(15 downto 0);
    signal conv131_383 : std_logic_vector(15 downto 0);
    signal conv134_396 : std_logic_vector(15 downto 0);
    signal conv144_483 : std_logic_vector(63 downto 0);
    signal conv149_496 : std_logic_vector(63 downto 0);
    signal conv155_514 : std_logic_vector(63 downto 0);
    signal conv161_532 : std_logic_vector(63 downto 0);
    signal conv167_550 : std_logic_vector(63 downto 0);
    signal conv173_568 : std_logic_vector(63 downto 0);
    signal conv179_586 : std_logic_vector(63 downto 0);
    signal conv17_82 : std_logic_vector(15 downto 0);
    signal conv185_604 : std_logic_vector(63 downto 0);
    signal conv1_32 : std_logic_vector(15 downto 0);
    signal conv200_690 : std_logic_vector(63 downto 0);
    signal conv205_703 : std_logic_vector(63 downto 0);
    signal conv20_95 : std_logic_vector(15 downto 0);
    signal conv211_721 : std_logic_vector(63 downto 0);
    signal conv217_739 : std_logic_vector(63 downto 0);
    signal conv223_757 : std_logic_vector(63 downto 0);
    signal conv229_775 : std_logic_vector(63 downto 0);
    signal conv235_793 : std_logic_vector(63 downto 0);
    signal conv241_811 : std_logic_vector(63 downto 0);
    signal conv253_844 : std_logic_vector(31 downto 0);
    signal conv255_848 : std_logic_vector(31 downto 0);
    signal conv258_852 : std_logic_vector(31 downto 0);
    signal conv26_107 : std_logic_vector(15 downto 0);
    signal conv29_120 : std_logic_vector(15 downto 0);
    signal conv302_1043 : std_logic_vector(15 downto 0);
    signal conv304_1050 : std_logic_vector(15 downto 0);
    signal conv319_1099 : std_logic_vector(15 downto 0);
    signal conv321_1106 : std_logic_vector(15 downto 0);
    signal conv336_1155 : std_logic_vector(15 downto 0);
    signal conv338_1162 : std_logic_vector(15 downto 0);
    signal conv35_132 : std_logic_vector(15 downto 0);
    signal conv365_1263 : std_logic_vector(7 downto 0);
    signal conv371_1273 : std_logic_vector(7 downto 0);
    signal conv377_1283 : std_logic_vector(7 downto 0);
    signal conv383_1293 : std_logic_vector(7 downto 0);
    signal conv389_1303 : std_logic_vector(7 downto 0);
    signal conv38_145 : std_logic_vector(15 downto 0);
    signal conv395_1313 : std_logic_vector(7 downto 0);
    signal conv3_45 : std_logic_vector(15 downto 0);
    signal conv401_1323 : std_logic_vector(7 downto 0);
    signal conv407_1333 : std_logic_vector(7 downto 0);
    signal conv44_157 : std_logic_vector(15 downto 0);
    signal conv47_170 : std_logic_vector(15 downto 0);
    signal conv53_182 : std_logic_vector(15 downto 0);
    signal conv56_195 : std_logic_vector(15 downto 0);
    signal conv61_204 : std_logic_vector(31 downto 0);
    signal conv63_208 : std_logic_vector(31 downto 0);
    signal conv65_212 : std_logic_vector(31 downto 0);
    signal conv82_249 : std_logic_vector(31 downto 0);
    signal conv84_253 : std_logic_vector(31 downto 0);
    signal conv87_257 : std_logic_vector(31 downto 0);
    signal conv8_57 : std_logic_vector(15 downto 0);
    signal conv90_261 : std_logic_vector(31 downto 0);
    signal conv95_283 : std_logic_vector(15 downto 0);
    signal conv98_296 : std_logic_vector(15 downto 0);
    signal exitcond1_1368 : std_logic_vector(0 downto 0);
    signal exitcond2_831 : std_logic_vector(0 downto 0);
    signal exitcond3_624 : std_logic_vector(0 downto 0);
    signal exitcond_943 : std_logic_vector(0 downto 0);
    signal iNsTr_14_234 : std_logic_vector(31 downto 0);
    signal iNsTr_187_1225 : std_logic_vector(63 downto 0);
    signal iNsTr_26_446 : std_logic_vector(63 downto 0);
    signal iNsTr_39_653 : std_logic_vector(63 downto 0);
    signal iNsTr_53_897 : std_logic_vector(63 downto 0);
    signal indvar453_913 : std_logic_vector(63 downto 0);
    signal indvar467_669 : std_logic_vector(63 downto 0);
    signal indvar483_462 : std_logic_vector(63 downto 0);
    signal indvar_1241 : std_logic_vector(63 downto 0);
    signal indvarx_xnext454_938 : std_logic_vector(63 downto 0);
    signal indvarx_xnext468_826 : std_logic_vector(63 downto 0);
    signal indvarx_xnext484_619 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1363 : std_logic_vector(63 downto 0);
    signal mul256_857 : std_logic_vector(31 downto 0);
    signal mul259_862 : std_logic_vector(31 downto 0);
    signal mul66_222 : std_logic_vector(31 downto 0);
    signal mul85_266 : std_logic_vector(31 downto 0);
    signal mul88_271 : std_logic_vector(31 downto 0);
    signal mul91_276 : std_logic_vector(31 downto 0);
    signal mul_217 : std_logic_vector(31 downto 0);
    signal ptr_deref_1258_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1258_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1258_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1258_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1258_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_611_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_611_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_611_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_611_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_611_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_611_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_818_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_818_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_818_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_818_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_818_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_818_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_929_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_929_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_929_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_929_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_929_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_929_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_314 : std_logic_vector(15 downto 0);
    signal shl114_339 : std_logic_vector(15 downto 0);
    signal shl123_364 : std_logic_vector(15 downto 0);
    signal shl132_389 : std_logic_vector(15 downto 0);
    signal shl146_489 : std_logic_vector(63 downto 0);
    signal shl152_507 : std_logic_vector(63 downto 0);
    signal shl158_525 : std_logic_vector(63 downto 0);
    signal shl164_543 : std_logic_vector(63 downto 0);
    signal shl170_561 : std_logic_vector(63 downto 0);
    signal shl176_579 : std_logic_vector(63 downto 0);
    signal shl182_597 : std_logic_vector(63 downto 0);
    signal shl18_88 : std_logic_vector(15 downto 0);
    signal shl202_696 : std_logic_vector(63 downto 0);
    signal shl208_714 : std_logic_vector(63 downto 0);
    signal shl214_732 : std_logic_vector(63 downto 0);
    signal shl220_750 : std_logic_vector(63 downto 0);
    signal shl226_768 : std_logic_vector(63 downto 0);
    signal shl232_786 : std_logic_vector(63 downto 0);
    signal shl238_804 : std_logic_vector(63 downto 0);
    signal shl27_113 : std_logic_vector(15 downto 0);
    signal shl36_138 : std_logic_vector(15 downto 0);
    signal shl45_163 : std_logic_vector(15 downto 0);
    signal shl54_188 : std_logic_vector(15 downto 0);
    signal shl96_289 : std_logic_vector(15 downto 0);
    signal shl9_63 : std_logic_vector(15 downto 0);
    signal shl_38 : std_logic_vector(15 downto 0);
    signal shr301_1039 : std_logic_vector(31 downto 0);
    signal shr318_1095 : std_logic_vector(31 downto 0);
    signal shr335_1151 : std_logic_vector(31 downto 0);
    signal shr368_1269 : std_logic_vector(63 downto 0);
    signal shr374_1279 : std_logic_vector(63 downto 0);
    signal shr380_1289 : std_logic_vector(63 downto 0);
    signal shr386_1299 : std_logic_vector(63 downto 0);
    signal shr392_1309 : std_logic_vector(63 downto 0);
    signal shr398_1319 : std_logic_vector(63 downto 0);
    signal shr404_1329 : std_logic_vector(63 downto 0);
    signal shr_228 : std_logic_vector(31 downto 0);
    signal tmp362_1259 : std_logic_vector(63 downto 0);
    signal tmp448_1209 : std_logic_vector(31 downto 0);
    signal tmp448x_xop_1221 : std_logic_vector(31 downto 0);
    signal tmp449_1215 : std_logic_vector(0 downto 0);
    signal tmp452_1238 : std_logic_vector(63 downto 0);
    signal tmp460_881 : std_logic_vector(31 downto 0);
    signal tmp460x_xop_893 : std_logic_vector(31 downto 0);
    signal tmp461_887 : std_logic_vector(0 downto 0);
    signal tmp465_910 : std_logic_vector(63 downto 0);
    signal tmp476_637 : std_logic_vector(31 downto 0);
    signal tmp476x_xop_649 : std_logic_vector(31 downto 0);
    signal tmp477_643 : std_logic_vector(0 downto 0);
    signal tmp481_666 : std_logic_vector(63 downto 0);
    signal tmp490x_xop_442 : std_logic_vector(31 downto 0);
    signal tmp491_436 : std_logic_vector(0 downto 0);
    signal tmp495_459 : std_logic_vector(63 downto 0);
    signal type_cast_1037_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1093_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_111_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1149_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1190_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1194_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1207_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1213_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1219_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1229_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1247_wire : std_logic_vector(63 downto 0);
    signal type_cast_1267_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1277_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1287_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1297_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1307_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1317_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1327_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1361_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_136_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_161_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_186_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_226_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_232_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_238_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_287_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_312_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_337_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_362_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_36_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_387_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_405_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_421_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_434_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_440_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_450_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_466_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_468_wire : std_logic_vector(63 downto 0);
    signal type_cast_487_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_505_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_523_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_541_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_559_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_577_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_595_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_617_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_61_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_635_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_657_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_672_wire : std_logic_vector(63 downto 0);
    signal type_cast_675_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_694_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_712_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_730_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_748_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_766_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_784_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_802_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_866_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_86_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_879_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_885_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_901_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_916_wire : std_logic_vector(63 downto 0);
    signal type_cast_919_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_931_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_936_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_960_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_992_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_996_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop497_903 : std_logic_vector(63 downto 0);
    signal xx_xop498_659 : std_logic_vector(63 downto 0);
    signal xx_xop499_452 : std_logic_vector(63 downto 0);
    signal xx_xop_1231 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1253_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1253_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1253_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1253_resized_base_address <= "00000000000000";
    array_obj_ref_474_constant_part_of_offset <= "00000000000000";
    array_obj_ref_474_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_474_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_474_resized_base_address <= "00000000000000";
    array_obj_ref_681_constant_part_of_offset <= "00000100010";
    array_obj_ref_681_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_681_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_681_resized_base_address <= "00000000000";
    array_obj_ref_925_constant_part_of_offset <= "00000000000000";
    array_obj_ref_925_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_925_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_925_resized_base_address <= "00000000000000";
    ptr_deref_1258_word_offset_0 <= "00000000000000";
    ptr_deref_611_word_offset_0 <= "00000000000000";
    ptr_deref_818_word_offset_0 <= "00000000000";
    ptr_deref_929_word_offset_0 <= "00000000000000";
    type_cast_1037_wire_constant <= "00000000000000000000000000010010";
    type_cast_1093_wire_constant <= "00000000000000000000000000010001";
    type_cast_111_wire_constant <= "0000000000001000";
    type_cast_1149_wire_constant <= "00000000000000000000000000010000";
    type_cast_1190_wire_constant <= "11111111";
    type_cast_1194_wire_constant <= "11111111";
    type_cast_1207_wire_constant <= "00000000000000000000000000000010";
    type_cast_1213_wire_constant <= "00000000000000000000000000000001";
    type_cast_1219_wire_constant <= "11111111111111111111111111111111";
    type_cast_1229_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1236_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1267_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1277_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1287_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1297_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1307_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1317_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1327_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1361_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_136_wire_constant <= "0000000000001000";
    type_cast_161_wire_constant <= "0000000000001000";
    type_cast_186_wire_constant <= "0000000000001000";
    type_cast_226_wire_constant <= "00000000000000000000000000000010";
    type_cast_232_wire_constant <= "00000000000000000000000000000001";
    type_cast_238_wire_constant <= "01111111111111111111111111111110";
    type_cast_287_wire_constant <= "0000000000001000";
    type_cast_312_wire_constant <= "0000000000001000";
    type_cast_337_wire_constant <= "0000000000001000";
    type_cast_362_wire_constant <= "0000000000001000";
    type_cast_36_wire_constant <= "0000000000001000";
    type_cast_387_wire_constant <= "0000000000001000";
    type_cast_405_wire_constant <= "00000000000000000000000000000011";
    type_cast_421_wire_constant <= "00000000000000000000000000000011";
    type_cast_434_wire_constant <= "00000000000000000000000000000001";
    type_cast_440_wire_constant <= "11111111111111111111111111111111";
    type_cast_450_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_466_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_487_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_505_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_523_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_541_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_559_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_577_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_595_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_617_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_61_wire_constant <= "0000000000001000";
    type_cast_635_wire_constant <= "00000000000000000000000000000010";
    type_cast_641_wire_constant <= "00000000000000000000000000000001";
    type_cast_647_wire_constant <= "11111111111111111111111111111111";
    type_cast_657_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_664_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_675_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_694_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_712_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_730_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_748_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_766_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_784_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_802_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_824_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_866_wire_constant <= "00000000000000000000000000000011";
    type_cast_86_wire_constant <= "0000000000001000";
    type_cast_879_wire_constant <= "00000000000000000000000000000010";
    type_cast_885_wire_constant <= "00000000000000000000000000000001";
    type_cast_891_wire_constant <= "11111111111111111111111111111111";
    type_cast_901_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_919_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_931_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_936_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_956_wire_constant <= "11111111";
    type_cast_960_wire_constant <= "11111111";
    type_cast_992_wire_constant <= "0000000000000000";
    type_cast_996_wire_constant <= "0000000000000000";
    phi_stmt_1241: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1245_wire_constant & type_cast_1247_wire;
      req <= phi_stmt_1241_req_0 & phi_stmt_1241_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1241",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1241_ack_0,
          idata => idata,
          odata => indvar_1241,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1241
    phi_stmt_462: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_466_wire_constant & type_cast_468_wire;
      req <= phi_stmt_462_req_0 & phi_stmt_462_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_462",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_462_ack_0,
          idata => idata,
          odata => indvar483_462,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_462
    phi_stmt_669: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_672_wire & type_cast_675_wire_constant;
      req <= phi_stmt_669_req_0 & phi_stmt_669_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_669",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_669_ack_0,
          idata => idata,
          odata => indvar467_669,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_669
    phi_stmt_913: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_916_wire & type_cast_919_wire_constant;
      req <= phi_stmt_913_req_0 & phi_stmt_913_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_913",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_913_ack_0,
          idata => idata,
          odata => indvar453_913,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_913
    -- flow-through select operator MUX_1237_inst
    tmp452_1238 <= xx_xop_1231 when (tmp449_1215(0) /=  '0') else type_cast_1236_wire_constant;
    -- flow-through select operator MUX_458_inst
    tmp495_459 <= xx_xop499_452 when (tmp491_436(0) /=  '0') else type_cast_457_wire_constant;
    -- flow-through select operator MUX_665_inst
    tmp481_666 <= xx_xop498_659 when (tmp477_643(0) /=  '0') else type_cast_664_wire_constant;
    -- flow-through select operator MUX_909_inst
    tmp465_910 <= xx_xop497_903 when (tmp461_887(0) /=  '0') else type_cast_908_wire_constant;
    addr_of_1254_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1254_final_reg_req_0;
      addr_of_1254_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1254_final_reg_req_1;
      addr_of_1254_final_reg_ack_1<= rack(0);
      addr_of_1254_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1254_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1253_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx361_1255,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_475_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_475_final_reg_req_0;
      addr_of_475_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_475_final_reg_req_1;
      addr_of_475_final_reg_ack_1<= rack(0);
      addr_of_475_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_475_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_474_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_476,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_682_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_682_final_reg_req_0;
      addr_of_682_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_682_final_reg_req_1;
      addr_of_682_final_reg_ack_1<= rack(0);
      addr_of_682_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_682_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_681_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_683,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_926_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_926_final_reg_req_0;
      addr_of_926_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_926_final_reg_req_1;
      addr_of_926_final_reg_ack_1<= rack(0);
      addr_of_926_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_926_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_925_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1042_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1042_inst_req_0;
      type_cast_1042_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1042_inst_req_1;
      type_cast_1042_inst_ack_1<= rack(0);
      type_cast_1042_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1042_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr301_1039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv302_1043,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1049_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1049_inst_req_0;
      type_cast_1049_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1049_inst_req_1;
      type_cast_1049_inst_ack_1<= rack(0);
      type_cast_1049_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1049_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_1050,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_106_inst_req_0;
      type_cast_106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_106_inst_req_1;
      type_cast_106_inst_ack_1<= rack(0);
      type_cast_106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1098_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1098_inst_req_0;
      type_cast_1098_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1098_inst_req_1;
      type_cast_1098_inst_ack_1<= rack(0);
      type_cast_1098_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1098_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr318_1095,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv319_1099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1105_inst_req_0;
      type_cast_1105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1105_inst_req_1;
      type_cast_1105_inst_ack_1<= rack(0);
      type_cast_1105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv321_1106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1154_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1154_inst_req_0;
      type_cast_1154_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1154_inst_req_1;
      type_cast_1154_inst_ack_1<= rack(0);
      type_cast_1154_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1154_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr335_1151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv336_1155,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1161_inst_req_0;
      type_cast_1161_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1161_inst_req_1;
      type_cast_1161_inst_ack_1<= rack(0);
      type_cast_1161_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv338_1162,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_119_inst_req_0;
      type_cast_119_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_119_inst_req_1;
      type_cast_119_inst_ack_1<= rack(0);
      type_cast_119_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_116,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1224_inst_req_0;
      type_cast_1224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1224_inst_req_1;
      type_cast_1224_inst_ack_1<= rack(0);
      type_cast_1224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp448x_xop_1221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_187_1225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1247_inst_req_0;
      type_cast_1247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1247_inst_req_1;
      type_cast_1247_inst_ack_1<= rack(0);
      type_cast_1247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1247_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1262_inst_req_0;
      type_cast_1262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1262_inst_req_1;
      type_cast_1262_inst_ack_1<= rack(0);
      type_cast_1262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp362_1259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv365_1263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1272_inst_req_0;
      type_cast_1272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1272_inst_req_1;
      type_cast_1272_inst_ack_1<= rack(0);
      type_cast_1272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr368_1269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv371_1273,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1282_inst_req_0;
      type_cast_1282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1282_inst_req_1;
      type_cast_1282_inst_ack_1<= rack(0);
      type_cast_1282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr374_1279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv377_1283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1292_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1292_inst_req_0;
      type_cast_1292_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1292_inst_req_1;
      type_cast_1292_inst_ack_1<= rack(0);
      type_cast_1292_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1292_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr380_1289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv383_1293,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1302_inst_req_0;
      type_cast_1302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1302_inst_req_1;
      type_cast_1302_inst_ack_1<= rack(0);
      type_cast_1302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr386_1299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv389_1303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1312_inst_req_0;
      type_cast_1312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1312_inst_req_1;
      type_cast_1312_inst_ack_1<= rack(0);
      type_cast_1312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr392_1309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv395_1313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_131_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_131_inst_req_0;
      type_cast_131_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_131_inst_req_1;
      type_cast_131_inst_ack_1<= rack(0);
      type_cast_131_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_131_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1322_inst_req_0;
      type_cast_1322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1322_inst_req_1;
      type_cast_1322_inst_ack_1<= rack(0);
      type_cast_1322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr398_1319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv401_1323,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1332_inst_req_0;
      type_cast_1332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1332_inst_req_1;
      type_cast_1332_inst_ack_1<= rack(0);
      type_cast_1332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr404_1329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv407_1333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_144_inst_req_0;
      type_cast_144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_144_inst_req_1;
      type_cast_144_inst_ack_1<= rack(0);
      type_cast_144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_156_inst_req_0;
      type_cast_156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_156_inst_req_1;
      type_cast_156_inst_ack_1<= rack(0);
      type_cast_156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_169_inst_req_0;
      type_cast_169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_169_inst_req_1;
      type_cast_169_inst_ack_1<= rack(0);
      type_cast_169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_166,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_181_inst_req_0;
      type_cast_181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_181_inst_req_1;
      type_cast_181_inst_ack_1<= rack(0);
      type_cast_181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_178,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_194_inst_req_0;
      type_cast_194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_194_inst_req_1;
      type_cast_194_inst_ack_1<= rack(0);
      type_cast_194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_203_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_203_inst_req_0;
      type_cast_203_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_203_inst_req_1;
      type_cast_203_inst_ack_1<= rack(0);
      type_cast_203_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_203_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_50,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_204,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_207_inst_req_0;
      type_cast_207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_207_inst_req_1;
      type_cast_207_inst_ack_1<= rack(0);
      type_cast_207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_75,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_248_inst_req_0;
      type_cast_248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_248_inst_req_1;
      type_cast_248_inst_ack_1<= rack(0);
      type_cast_248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_249,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_252_inst_req_0;
      type_cast_252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_252_inst_req_1;
      type_cast_252_inst_ack_1<= rack(0);
      type_cast_252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_150,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_256_inst_req_0;
      type_cast_256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_256_inst_req_1;
      type_cast_256_inst_ack_1<= rack(0);
      type_cast_256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_260_inst_req_0;
      type_cast_260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_260_inst_req_1;
      type_cast_260_inst_ack_1<= rack(0);
      type_cast_260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_282_inst_req_0;
      type_cast_282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_282_inst_req_1;
      type_cast_282_inst_ack_1<= rack(0);
      type_cast_282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_295_inst_req_0;
      type_cast_295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_295_inst_req_1;
      type_cast_295_inst_ack_1<= rack(0);
      type_cast_295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_307_inst_req_0;
      type_cast_307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_307_inst_req_1;
      type_cast_307_inst_ack_1<= rack(0);
      type_cast_307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_307_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_308,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_31_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_31_inst_req_0;
      type_cast_31_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_31_inst_req_1;
      type_cast_31_inst_ack_1<= rack(0);
      type_cast_31_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_31_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_28,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_32,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_320_inst_req_0;
      type_cast_320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_320_inst_req_1;
      type_cast_320_inst_ack_1<= rack(0);
      type_cast_320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_332_inst_req_0;
      type_cast_332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_332_inst_req_1;
      type_cast_332_inst_ack_1<= rack(0);
      type_cast_332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_382_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_382_inst_req_0;
      type_cast_382_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_382_inst_req_1;
      type_cast_382_inst_ack_1<= rack(0);
      type_cast_382_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_382_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_379,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_383,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_395_inst_req_0;
      type_cast_395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_395_inst_req_1;
      type_cast_395_inst_ack_1<= rack(0);
      type_cast_395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_445_inst_req_0;
      type_cast_445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_445_inst_req_1;
      type_cast_445_inst_ack_1<= rack(0);
      type_cast_445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp490x_xop_442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_44_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_44_inst_req_0;
      type_cast_44_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_44_inst_req_1;
      type_cast_44_inst_ack_1<= rack(0);
      type_cast_44_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_44_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_45,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_468_inst_req_0;
      type_cast_468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_468_inst_req_1;
      type_cast_468_inst_ack_1<= rack(0);
      type_cast_468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_468_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext484_619,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_468_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_482_inst_req_0;
      type_cast_482_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_482_inst_req_1;
      type_cast_482_inst_ack_1<= rack(0);
      type_cast_482_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_482_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_479,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_495_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_495_inst_req_0;
      type_cast_495_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_495_inst_req_1;
      type_cast_495_inst_ack_1<= rack(0);
      type_cast_495_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_495_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_496,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_513_inst_req_0;
      type_cast_513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_513_inst_req_1;
      type_cast_513_inst_ack_1<= rack(0);
      type_cast_513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_510,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_531_inst_req_0;
      type_cast_531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_531_inst_req_1;
      type_cast_531_inst_ack_1<= rack(0);
      type_cast_531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_528,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_549_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_549_inst_req_0;
      type_cast_549_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_549_inst_req_1;
      type_cast_549_inst_ack_1<= rack(0);
      type_cast_549_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_549_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_546,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_550,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_567_inst_req_0;
      type_cast_567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_567_inst_req_1;
      type_cast_567_inst_ack_1<= rack(0);
      type_cast_567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_564,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_568,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_56_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_56_inst_req_0;
      type_cast_56_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_56_inst_req_1;
      type_cast_56_inst_ack_1<= rack(0);
      type_cast_56_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_56_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_53,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_57,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_585_inst_req_0;
      type_cast_585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_585_inst_req_1;
      type_cast_585_inst_ack_1<= rack(0);
      type_cast_585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_582,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_603_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_603_inst_req_0;
      type_cast_603_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_603_inst_req_1;
      type_cast_603_inst_ack_1<= rack(0);
      type_cast_603_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_603_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_600,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_604,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_652_inst_req_0;
      type_cast_652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_652_inst_req_1;
      type_cast_652_inst_ack_1<= rack(0);
      type_cast_652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp476x_xop_649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_672_inst_req_0;
      type_cast_672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_672_inst_req_1;
      type_cast_672_inst_ack_1<= rack(0);
      type_cast_672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext468_826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_672_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_689_inst_req_0;
      type_cast_689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_689_inst_req_1;
      type_cast_689_inst_ack_1<= rack(0);
      type_cast_689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_69_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_69_inst_req_0;
      type_cast_69_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_69_inst_req_1;
      type_cast_69_inst_ack_1<= rack(0);
      type_cast_69_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_69_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_66,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_70,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_702_inst_req_0;
      type_cast_702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_702_inst_req_1;
      type_cast_702_inst_ack_1<= rack(0);
      type_cast_702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_703,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_720_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_720_inst_req_0;
      type_cast_720_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_720_inst_req_1;
      type_cast_720_inst_ack_1<= rack(0);
      type_cast_720_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_720_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_717,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_721,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_738_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_738_inst_req_0;
      type_cast_738_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_738_inst_req_1;
      type_cast_738_inst_ack_1<= rack(0);
      type_cast_738_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_738_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_739,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_756_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_756_inst_req_0;
      type_cast_756_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_756_inst_req_1;
      type_cast_756_inst_ack_1<= rack(0);
      type_cast_756_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_756_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_753,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_774_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_774_inst_req_0;
      type_cast_774_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_774_inst_req_1;
      type_cast_774_inst_ack_1<= rack(0);
      type_cast_774_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_774_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_771,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_775,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_792_inst_req_0;
      type_cast_792_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_792_inst_req_1;
      type_cast_792_inst_ack_1<= rack(0);
      type_cast_792_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_792_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_793,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_810_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_810_inst_req_0;
      type_cast_810_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_810_inst_req_1;
      type_cast_810_inst_ack_1<= rack(0);
      type_cast_810_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_810_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_811,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_81_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_81_inst_req_0;
      type_cast_81_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_81_inst_req_1;
      type_cast_81_inst_ack_1<= rack(0);
      type_cast_81_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_81_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_78,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_82,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_843_inst_req_0;
      type_cast_843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_843_inst_req_1;
      type_cast_843_inst_ack_1<= rack(0);
      type_cast_843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_351,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_847_inst_req_0;
      type_cast_847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_847_inst_req_1;
      type_cast_847_inst_ack_1<= rack(0);
      type_cast_847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_847_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_401,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_896_inst_req_0;
      type_cast_896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_896_inst_req_1;
      type_cast_896_inst_ack_1<= rack(0);
      type_cast_896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp460x_xop_893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_897,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_916_inst_req_0;
      type_cast_916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_916_inst_req_1;
      type_cast_916_inst_ack_1<= rack(0);
      type_cast_916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext454_938,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_916_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_94_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_94_inst_req_0;
      type_cast_94_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_94_inst_req_1;
      type_cast_94_inst_ack_1<= rack(0);
      type_cast_94_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_94_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_91,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1253_index_1_rename
    process(R_indvar_1252_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1252_resized;
      ov(13 downto 0) := iv;
      R_indvar_1252_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1253_index_1_resize
    process(indvar_1241) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1241;
      ov := iv(13 downto 0);
      R_indvar_1252_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1253_root_address_inst
    process(array_obj_ref_1253_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1253_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1253_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_474_index_1_rename
    process(R_indvar483_473_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar483_473_resized;
      ov(13 downto 0) := iv;
      R_indvar483_473_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_474_index_1_resize
    process(indvar483_462) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar483_462;
      ov := iv(13 downto 0);
      R_indvar483_473_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_474_root_address_inst
    process(array_obj_ref_474_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_474_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_474_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_681_index_1_rename
    process(R_indvar467_680_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar467_680_resized;
      ov(10 downto 0) := iv;
      R_indvar467_680_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_681_index_1_resize
    process(indvar467_669) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar467_669;
      ov := iv(10 downto 0);
      R_indvar467_680_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_681_root_address_inst
    process(array_obj_ref_681_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_681_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_681_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_925_index_1_rename
    process(R_indvar453_924_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar453_924_resized;
      ov(13 downto 0) := iv;
      R_indvar453_924_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_925_index_1_resize
    process(indvar453_913) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar453_913;
      ov := iv(13 downto 0);
      R_indvar453_924_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_925_root_address_inst
    process(array_obj_ref_925_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_925_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_925_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1258_addr_0
    process(ptr_deref_1258_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1258_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1258_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1258_base_resize
    process(arrayidx361_1255) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx361_1255;
      ov := iv(13 downto 0);
      ptr_deref_1258_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1258_gather_scatter
    process(ptr_deref_1258_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1258_data_0;
      ov(63 downto 0) := iv;
      tmp362_1259 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1258_root_address_inst
    process(ptr_deref_1258_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1258_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1258_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_611_addr_0
    process(ptr_deref_611_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_611_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_611_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_611_base_resize
    process(arrayidx_476) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_476;
      ov := iv(13 downto 0);
      ptr_deref_611_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_611_gather_scatter
    process(add186_609) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_609;
      ov(63 downto 0) := iv;
      ptr_deref_611_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_611_root_address_inst
    process(ptr_deref_611_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_611_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_611_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_818_addr_0
    process(ptr_deref_818_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_818_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_818_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_818_base_resize
    process(arrayidx246_683) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_683;
      ov := iv(10 downto 0);
      ptr_deref_818_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_818_gather_scatter
    process(add242_816) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_816;
      ov(63 downto 0) := iv;
      ptr_deref_818_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_818_root_address_inst
    process(ptr_deref_818_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_818_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_818_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_addr_0
    process(ptr_deref_929_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_929_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_929_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_base_resize
    process(arrayidx269_927) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_927;
      ov := iv(13 downto 0);
      ptr_deref_929_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_gather_scatter
    process(type_cast_931_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_931_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_929_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_root_address_inst
    process(ptr_deref_929_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_929_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_929_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1197_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264433_868;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1197_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1197_branch_req_0,
          ack0 => if_stmt_1197_branch_ack_0,
          ack1 => if_stmt_1197_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1369_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1368;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1369_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1369_branch_req_0,
          ack0 => if_stmt_1369_branch_ack_0,
          ack1 => if_stmt_1369_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_409_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp441_408;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_409_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_409_branch_req_0,
          ack0 => if_stmt_409_branch_ack_0,
          ack1 => if_stmt_409_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_424_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194437_423;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_424_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_424_branch_req_0,
          ack0 => if_stmt_424_branch_ack_0,
          ack1 => if_stmt_424_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_625_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_624;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_625_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_625_branch_req_0,
          ack0 => if_stmt_625_branch_ack_0,
          ack1 => if_stmt_625_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_832_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_831;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_832_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_832_branch_req_0,
          ack0 => if_stmt_832_branch_ack_0,
          ack1 => if_stmt_832_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_869_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264433_868;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_869_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_869_branch_req_0,
          ack0 => if_stmt_869_branch_ack_0,
          ack1 => if_stmt_869_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_944_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_943;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_944_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_944_branch_req_0,
          ack0 => if_stmt_944_branch_ack_0,
          ack1 => if_stmt_944_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1220_inst
    process(tmp448_1209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp448_1209, type_cast_1219_wire_constant, tmp_var);
      tmp448x_xop_1221 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_244_inst
    process(add74_240, shr_228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_240, shr_228, tmp_var);
      add79_245 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_441_inst
    process(shr_228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_228, type_cast_440_wire_constant, tmp_var);
      tmp490x_xop_442 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_648_inst
    process(tmp476_637) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp476_637, type_cast_647_wire_constant, tmp_var);
      tmp476x_xop_649 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_892_inst
    process(tmp460_881) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp460_881, type_cast_891_wire_constant, tmp_var);
      tmp460x_xop_893 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1230_inst
    process(iNsTr_187_1225) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_187_1225, type_cast_1229_wire_constant, tmp_var);
      xx_xop_1231 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1362_inst
    process(indvar_1241) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1241, type_cast_1361_wire_constant, tmp_var);
      indvarx_xnext_1363 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_451_inst
    process(iNsTr_26_446) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_446, type_cast_450_wire_constant, tmp_var);
      xx_xop499_452 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_618_inst
    process(indvar483_462) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar483_462, type_cast_617_wire_constant, tmp_var);
      indvarx_xnext484_619 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_658_inst
    process(iNsTr_39_653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_653, type_cast_657_wire_constant, tmp_var);
      xx_xop498_659 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_825_inst
    process(indvar467_669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar467_669, type_cast_824_wire_constant, tmp_var);
      indvarx_xnext468_826 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_902_inst
    process(iNsTr_53_897) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_897, type_cast_901_wire_constant, tmp_var);
      xx_xop497_903 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_937_inst
    process(indvar453_913) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar453_913, type_cast_936_wire_constant, tmp_var);
      indvarx_xnext454_938 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_239_inst
    process(iNsTr_14_234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_234, type_cast_238_wire_constant, tmp_var);
      add74_240 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1367_inst
    process(indvarx_xnext_1363, tmp452_1238) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1363, tmp452_1238, tmp_var);
      exitcond1_1368 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_623_inst
    process(indvarx_xnext484_619, tmp495_459) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext484_619, tmp495_459, tmp_var);
      exitcond3_624 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_830_inst
    process(indvarx_xnext468_826, tmp481_666) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext468_826, tmp481_666, tmp_var);
      exitcond2_831 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_942_inst
    process(indvarx_xnext454_938, tmp465_910) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext454_938, tmp465_910, tmp_var);
      exitcond_943 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1038_inst
    process(mul66_222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_222, type_cast_1037_wire_constant, tmp_var);
      shr301_1039 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1094_inst
    process(mul66_222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_222, type_cast_1093_wire_constant, tmp_var);
      shr318_1095 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1150_inst
    process(add79_245) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_245, type_cast_1149_wire_constant, tmp_var);
      shr335_1151 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1208_inst
    process(mul259_862) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_862, type_cast_1207_wire_constant, tmp_var);
      tmp448_1209 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_227_inst
    process(mul66_222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_222, type_cast_226_wire_constant, tmp_var);
      shr_228 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_233_inst
    process(mul66_222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_222, type_cast_232_wire_constant, tmp_var);
      iNsTr_14_234 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_636_inst
    process(mul91_276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_276, type_cast_635_wire_constant, tmp_var);
      tmp476_637 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_880_inst
    process(mul259_862) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_862, type_cast_879_wire_constant, tmp_var);
      tmp460_881 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1268_inst
    process(tmp362_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_1259, type_cast_1267_wire_constant, tmp_var);
      shr368_1269 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1278_inst
    process(tmp362_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_1259, type_cast_1277_wire_constant, tmp_var);
      shr374_1279 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1288_inst
    process(tmp362_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_1259, type_cast_1287_wire_constant, tmp_var);
      shr380_1289 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1298_inst
    process(tmp362_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_1259, type_cast_1297_wire_constant, tmp_var);
      shr386_1299 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1308_inst
    process(tmp362_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_1259, type_cast_1307_wire_constant, tmp_var);
      shr392_1309 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1318_inst
    process(tmp362_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_1259, type_cast_1317_wire_constant, tmp_var);
      shr398_1319 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1328_inst
    process(tmp362_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_1259, type_cast_1327_wire_constant, tmp_var);
      shr404_1329 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_216_inst
    process(conv63_208, conv61_204) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_208, conv61_204, tmp_var);
      mul_217 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_221_inst
    process(mul_217, conv65_212) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_217, conv65_212, tmp_var);
      mul66_222 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_265_inst
    process(conv84_253, conv82_249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_253, conv82_249, tmp_var);
      mul85_266 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_270_inst
    process(mul85_266, conv87_257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_266, conv87_257, tmp_var);
      mul88_271 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_275_inst
    process(mul88_271, conv90_261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_271, conv90_261, tmp_var);
      mul91_276 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_856_inst
    process(conv255_848, conv253_844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_848, conv253_844, tmp_var);
      mul256_857 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_861_inst
    process(mul256_857, conv258_852) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_857, conv258_852, tmp_var);
      mul259_862 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_124_inst
    process(shl27_113, conv29_120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_113, conv29_120, tmp_var);
      add30_125 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_149_inst
    process(shl36_138, conv38_145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_138, conv38_145, tmp_var);
      add39_150 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_174_inst
    process(shl45_163, conv47_170) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_163, conv47_170, tmp_var);
      add48_175 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_199_inst
    process(shl54_188, conv56_195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_188, conv56_195, tmp_var);
      add57_200 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_300_inst
    process(shl96_289, conv98_296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_289, conv98_296, tmp_var);
      add99_301 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_325_inst
    process(shl105_314, conv107_321) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_314, conv107_321, tmp_var);
      add108_326 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_350_inst
    process(shl114_339, conv116_346) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_339, conv116_346, tmp_var);
      add117_351 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_375_inst
    process(shl123_364, conv125_371) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_364, conv125_371, tmp_var);
      add126_376 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_400_inst
    process(shl132_389, conv134_396) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_389, conv134_396, tmp_var);
      add135_401 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_49_inst
    process(shl_38, conv3_45) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_38, conv3_45, tmp_var);
      add_50 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_74_inst
    process(shl9_63, conv11_70) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_63, conv11_70, tmp_var);
      add12_75 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_99_inst
    process(shl18_88, conv20_95) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_88, conv20_95, tmp_var);
      add21_100 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_500_inst
    process(shl146_489, conv149_496) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_489, conv149_496, tmp_var);
      add150_501 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_518_inst
    process(shl152_507, conv155_514) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_507, conv155_514, tmp_var);
      add156_519 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_536_inst
    process(shl158_525, conv161_532) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_525, conv161_532, tmp_var);
      add162_537 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_554_inst
    process(shl164_543, conv167_550) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_543, conv167_550, tmp_var);
      add168_555 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_572_inst
    process(shl170_561, conv173_568) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_561, conv173_568, tmp_var);
      add174_573 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_590_inst
    process(shl176_579, conv179_586) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_579, conv179_586, tmp_var);
      add180_591 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_608_inst
    process(shl182_597, conv185_604) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_597, conv185_604, tmp_var);
      add186_609 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_707_inst
    process(shl202_696, conv205_703) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_696, conv205_703, tmp_var);
      add206_708 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_725_inst
    process(shl208_714, conv211_721) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_714, conv211_721, tmp_var);
      add212_726 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_743_inst
    process(shl214_732, conv217_739) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_732, conv217_739, tmp_var);
      add218_744 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_761_inst
    process(shl220_750, conv223_757) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_750, conv223_757, tmp_var);
      add224_762 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_779_inst
    process(shl226_768, conv229_775) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_768, conv229_775, tmp_var);
      add230_780 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_797_inst
    process(shl232_786, conv235_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_786, conv235_793, tmp_var);
      add236_798 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_815_inst
    process(shl238_804, conv241_811) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_804, conv241_811, tmp_var);
      add242_816 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_112_inst
    process(conv26_107) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_107, type_cast_111_wire_constant, tmp_var);
      shl27_113 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_137_inst
    process(conv35_132) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_132, type_cast_136_wire_constant, tmp_var);
      shl36_138 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_162_inst
    process(conv44_157) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_157, type_cast_161_wire_constant, tmp_var);
      shl45_163 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_187_inst
    process(conv53_182) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_182, type_cast_186_wire_constant, tmp_var);
      shl54_188 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_288_inst
    process(conv95_283) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_283, type_cast_287_wire_constant, tmp_var);
      shl96_289 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_313_inst
    process(conv104_308) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_308, type_cast_312_wire_constant, tmp_var);
      shl105_314 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_338_inst
    process(conv113_333) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_333, type_cast_337_wire_constant, tmp_var);
      shl114_339 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_363_inst
    process(conv122_358) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_358, type_cast_362_wire_constant, tmp_var);
      shl123_364 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_37_inst
    process(conv1_32) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_32, type_cast_36_wire_constant, tmp_var);
      shl_38 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_388_inst
    process(conv131_383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_383, type_cast_387_wire_constant, tmp_var);
      shl132_389 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_62_inst
    process(conv8_57) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_57, type_cast_61_wire_constant, tmp_var);
      shl9_63 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_87_inst
    process(conv17_82) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_82, type_cast_86_wire_constant, tmp_var);
      shl18_88 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_488_inst
    process(conv144_483) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_483, type_cast_487_wire_constant, tmp_var);
      shl146_489 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_506_inst
    process(add150_501) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_501, type_cast_505_wire_constant, tmp_var);
      shl152_507 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_524_inst
    process(add156_519) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_519, type_cast_523_wire_constant, tmp_var);
      shl158_525 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_542_inst
    process(add162_537) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_537, type_cast_541_wire_constant, tmp_var);
      shl164_543 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_560_inst
    process(add168_555) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_555, type_cast_559_wire_constant, tmp_var);
      shl170_561 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_578_inst
    process(add174_573) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_573, type_cast_577_wire_constant, tmp_var);
      shl176_579 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_596_inst
    process(add180_591) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_591, type_cast_595_wire_constant, tmp_var);
      shl182_597 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_695_inst
    process(conv200_690) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_690, type_cast_694_wire_constant, tmp_var);
      shl202_696 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_713_inst
    process(add206_708) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_708, type_cast_712_wire_constant, tmp_var);
      shl208_714 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_731_inst
    process(add212_726) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_726, type_cast_730_wire_constant, tmp_var);
      shl214_732 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_749_inst
    process(add218_744) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_744, type_cast_748_wire_constant, tmp_var);
      shl220_750 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_767_inst
    process(add224_762) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_762, type_cast_766_wire_constant, tmp_var);
      shl226_768 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_785_inst
    process(add230_780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_780, type_cast_784_wire_constant, tmp_var);
      shl232_786 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_803_inst
    process(add236_798) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_798, type_cast_802_wire_constant, tmp_var);
      shl238_804 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1214_inst
    process(tmp448_1209) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp448_1209, type_cast_1213_wire_constant, tmp_var);
      tmp449_1215 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_406_inst
    process(mul66_222) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_222, type_cast_405_wire_constant, tmp_var);
      cmp441_408 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_422_inst
    process(mul91_276) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_276, type_cast_421_wire_constant, tmp_var);
      cmp194437_423 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_435_inst
    process(shr_228) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_228, type_cast_434_wire_constant, tmp_var);
      tmp491_436 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_642_inst
    process(tmp476_637) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp476_637, type_cast_641_wire_constant, tmp_var);
      tmp477_643 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_867_inst
    process(mul259_862) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_862, type_cast_866_wire_constant, tmp_var);
      cmp264433_868 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_886_inst
    process(tmp460_881) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp460_881, type_cast_885_wire_constant, tmp_var);
      tmp461_887 <= tmp_var; --
    end process;
    -- shared split operator group (99) : array_obj_ref_1253_index_offset 
    ApIntAdd_group_99: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1252_scaled;
      array_obj_ref_1253_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1253_index_offset_req_0;
      array_obj_ref_1253_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1253_index_offset_req_1;
      array_obj_ref_1253_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_99_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_99_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_99",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 99
    -- shared split operator group (100) : array_obj_ref_474_index_offset 
    ApIntAdd_group_100: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar483_473_scaled;
      array_obj_ref_474_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_474_index_offset_req_0;
      array_obj_ref_474_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_474_index_offset_req_1;
      array_obj_ref_474_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_100_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_100_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_100",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 100
    -- shared split operator group (101) : array_obj_ref_681_index_offset 
    ApIntAdd_group_101: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar467_680_scaled;
      array_obj_ref_681_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_681_index_offset_req_0;
      array_obj_ref_681_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_681_index_offset_req_1;
      array_obj_ref_681_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_101_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_101_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_101",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 101
    -- shared split operator group (102) : array_obj_ref_925_index_offset 
    ApIntAdd_group_102: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar453_924_scaled;
      array_obj_ref_925_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_925_index_offset_req_0;
      array_obj_ref_925_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_925_index_offset_req_1;
      array_obj_ref_925_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_102_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_102_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_102",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared load operator group (0) : ptr_deref_1258_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1258_load_0_req_0;
      ptr_deref_1258_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1258_load_0_req_1;
      ptr_deref_1258_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1258_word_address_0;
      ptr_deref_1258_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_611_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_611_store_0_req_0;
      ptr_deref_611_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_611_store_0_req_1;
      ptr_deref_611_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_611_word_address_0;
      data_in <= ptr_deref_611_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_818_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_818_store_0_req_0;
      ptr_deref_818_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_818_store_0_req_1;
      ptr_deref_818_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_818_word_address_0;
      data_in <= ptr_deref_818_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(10 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_929_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_929_store_0_req_0;
      ptr_deref_929_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_929_store_0_req_1;
      ptr_deref_929_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_929_word_address_0;
      data_in <= ptr_deref_929_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1176_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1176_inst_req_0;
      RPIPE_Block0_done_1176_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1176_inst_req_1;
      RPIPE_Block0_done_1176_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call343_1177 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1179_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1179_inst_req_0;
      RPIPE_Block1_done_1179_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1179_inst_req_1;
      RPIPE_Block1_done_1179_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call345_1180 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1182_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1182_inst_req_0;
      RPIPE_Block2_done_1182_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1182_inst_req_1;
      RPIPE_Block2_done_1182_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call347_1183 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1185_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1185_inst_req_0;
      RPIPE_Block3_done_1185_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1185_inst_req_1;
      RPIPE_Block3_done_1185_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call349_1186 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_102_inst RPIPE_ConvTranspose_input_pipe_152_inst RPIPE_ConvTranspose_input_pipe_190_inst RPIPE_ConvTranspose_input_pipe_52_inst RPIPE_ConvTranspose_input_pipe_115_inst RPIPE_ConvTranspose_input_pipe_177_inst RPIPE_ConvTranspose_input_pipe_65_inst RPIPE_ConvTranspose_input_pipe_77_inst RPIPE_ConvTranspose_input_pipe_127_inst RPIPE_ConvTranspose_input_pipe_90_inst RPIPE_ConvTranspose_input_pipe_140_inst RPIPE_ConvTranspose_input_pipe_40_inst RPIPE_ConvTranspose_input_pipe_27_inst RPIPE_ConvTranspose_input_pipe_165_inst RPIPE_ConvTranspose_input_pipe_491_inst RPIPE_ConvTranspose_input_pipe_545_inst RPIPE_ConvTranspose_input_pipe_478_inst RPIPE_ConvTranspose_input_pipe_563_inst RPIPE_ConvTranspose_input_pipe_366_inst RPIPE_ConvTranspose_input_pipe_509_inst RPIPE_ConvTranspose_input_pipe_527_inst RPIPE_ConvTranspose_input_pipe_378_inst RPIPE_ConvTranspose_input_pipe_391_inst RPIPE_ConvTranspose_input_pipe_353_inst RPIPE_ConvTranspose_input_pipe_341_inst RPIPE_ConvTranspose_input_pipe_328_inst RPIPE_ConvTranspose_input_pipe_316_inst RPIPE_ConvTranspose_input_pipe_303_inst RPIPE_ConvTranspose_input_pipe_291_inst RPIPE_ConvTranspose_input_pipe_278_inst RPIPE_ConvTranspose_input_pipe_581_inst RPIPE_ConvTranspose_input_pipe_599_inst RPIPE_ConvTranspose_input_pipe_685_inst RPIPE_ConvTranspose_input_pipe_698_inst RPIPE_ConvTranspose_input_pipe_716_inst RPIPE_ConvTranspose_input_pipe_734_inst RPIPE_ConvTranspose_input_pipe_752_inst RPIPE_ConvTranspose_input_pipe_770_inst RPIPE_ConvTranspose_input_pipe_788_inst RPIPE_ConvTranspose_input_pipe_806_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_102_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_152_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_52_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_177_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_77_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_127_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_27_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_491_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_545_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_478_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_563_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_509_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_527_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_378_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_353_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_328_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_303_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_278_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_581_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_599_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_685_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_698_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_716_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_734_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_752_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_770_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_788_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_806_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_102_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_152_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_52_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_177_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_77_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_127_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_27_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_491_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_545_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_478_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_563_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_509_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_527_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_378_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_353_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_328_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_303_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_278_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_581_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_599_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_685_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_698_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_716_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_734_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_752_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_770_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_788_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_806_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_102_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_152_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_52_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_177_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_77_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_127_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_27_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_491_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_545_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_478_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_563_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_509_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_527_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_378_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_353_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_328_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_303_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_278_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_581_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_599_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_685_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_698_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_716_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_734_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_752_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_770_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_788_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_806_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_102_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_152_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_52_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_177_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_77_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_127_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_27_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_491_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_545_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_478_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_563_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_509_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_527_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_378_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_353_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_328_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_303_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_278_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_581_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_599_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_685_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_698_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_716_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_734_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_752_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_770_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_788_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_806_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call23_103 <= data_out(319 downto 312);
      call41_153 <= data_out(311 downto 304);
      call55_191 <= data_out(303 downto 296);
      call5_53 <= data_out(295 downto 288);
      call28_116 <= data_out(287 downto 280);
      call50_178 <= data_out(279 downto 272);
      call10_66 <= data_out(271 downto 264);
      call14_78 <= data_out(263 downto 256);
      call32_128 <= data_out(255 downto 248);
      call19_91 <= data_out(247 downto 240);
      call37_141 <= data_out(239 downto 232);
      call2_41 <= data_out(231 downto 224);
      call_28 <= data_out(223 downto 216);
      call46_166 <= data_out(215 downto 208);
      call147_492 <= data_out(207 downto 200);
      call165_546 <= data_out(199 downto 192);
      call143_479 <= data_out(191 downto 184);
      call171_564 <= data_out(183 downto 176);
      call124_367 <= data_out(175 downto 168);
      call153_510 <= data_out(167 downto 160);
      call159_528 <= data_out(159 downto 152);
      call128_379 <= data_out(151 downto 144);
      call133_392 <= data_out(143 downto 136);
      call119_354 <= data_out(135 downto 128);
      call115_342 <= data_out(127 downto 120);
      call110_329 <= data_out(119 downto 112);
      call106_317 <= data_out(111 downto 104);
      call101_304 <= data_out(103 downto 96);
      call97_292 <= data_out(95 downto 88);
      call92_279 <= data_out(87 downto 80);
      call177_582 <= data_out(79 downto 72);
      call183_600 <= data_out(71 downto 64);
      call199_686 <= data_out(63 downto 56);
      call203_699 <= data_out(55 downto 48);
      call209_717 <= data_out(47 downto 40);
      call215_735 <= data_out(39 downto 32);
      call221_753 <= data_out(31 downto 24);
      call227_771 <= data_out(23 downto 16);
      call233_789 <= data_out(15 downto 8);
      call239_807 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_963_inst WPIPE_Block0_start_966_inst WPIPE_Block0_start_969_inst WPIPE_Block0_start_972_inst WPIPE_Block0_start_975_inst WPIPE_Block0_start_978_inst WPIPE_Block0_start_981_inst WPIPE_Block0_start_984_inst WPIPE_Block0_start_987_inst WPIPE_Block0_start_990_inst WPIPE_Block0_start_994_inst WPIPE_Block0_start_998_inst WPIPE_Block0_start_1001_inst WPIPE_Block0_start_1004_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_963_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_966_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_969_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_972_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_975_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_978_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_981_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_984_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_987_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_990_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_994_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_998_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_1001_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_1004_inst_req_0;
      WPIPE_Block0_start_963_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_966_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_969_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_972_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_975_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_978_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_981_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_984_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_987_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_990_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_994_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_998_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_1001_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_1004_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_963_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_966_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_969_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_972_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_975_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_978_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_981_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_984_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_987_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_990_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_994_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_998_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_1001_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_1004_inst_req_1;
      WPIPE_Block0_start_963_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_966_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_969_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_972_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_975_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_978_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_981_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_984_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_987_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_990_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_994_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_998_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_1001_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_1004_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_50 & add12_75 & add21_100 & add30_125 & add39_150 & add48_175 & add57_200 & add99_301 & add108_326 & type_cast_992_wire_constant & type_cast_996_wire_constant & add117_351 & add126_376 & add135_401;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1007_inst WPIPE_Block1_start_1010_inst WPIPE_Block1_start_1013_inst WPIPE_Block1_start_1016_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1022_inst WPIPE_Block1_start_1025_inst WPIPE_Block1_start_1028_inst WPIPE_Block1_start_1031_inst WPIPE_Block1_start_1044_inst WPIPE_Block1_start_1051_inst WPIPE_Block1_start_1054_inst WPIPE_Block1_start_1057_inst WPIPE_Block1_start_1060_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1007_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1010_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1013_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1016_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1022_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1025_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1028_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1031_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1044_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1051_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1054_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1057_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1060_inst_req_0;
      WPIPE_Block1_start_1007_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1010_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1013_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1016_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1025_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1028_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1031_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1044_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1051_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1054_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1057_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1060_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1007_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1010_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1013_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1016_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1022_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1025_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1028_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1031_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1044_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1051_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1054_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1057_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1060_inst_req_1;
      WPIPE_Block1_start_1007_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1010_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1013_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1016_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1025_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1028_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1031_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1044_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1051_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1054_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1057_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1060_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_50 & add12_75 & add21_100 & add30_125 & add39_150 & add48_175 & add57_200 & add99_301 & add108_326 & conv302_1043 & conv304_1050 & add117_351 & add126_376 & add135_401;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1063_inst WPIPE_Block2_start_1066_inst WPIPE_Block2_start_1069_inst WPIPE_Block2_start_1072_inst WPIPE_Block2_start_1075_inst WPIPE_Block2_start_1078_inst WPIPE_Block2_start_1081_inst WPIPE_Block2_start_1084_inst WPIPE_Block2_start_1087_inst WPIPE_Block2_start_1100_inst WPIPE_Block2_start_1107_inst WPIPE_Block2_start_1110_inst WPIPE_Block2_start_1113_inst WPIPE_Block2_start_1116_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1063_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1066_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1069_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1072_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1075_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1078_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1081_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1084_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1087_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1100_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1107_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1110_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1113_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1116_inst_req_0;
      WPIPE_Block2_start_1063_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1066_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1069_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1072_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1075_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1078_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1081_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1084_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1087_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1100_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1107_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1110_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1113_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1116_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1063_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1066_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1069_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1072_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1075_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1078_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1081_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1084_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1087_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1100_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1107_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1110_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1113_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1116_inst_req_1;
      WPIPE_Block2_start_1063_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1066_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1069_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1072_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1075_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1078_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1081_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1084_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1087_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1100_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1107_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1110_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1113_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1116_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_50 & add12_75 & add21_100 & add30_125 & add39_150 & add48_175 & add57_200 & add99_301 & add108_326 & conv319_1099 & conv321_1106 & add117_351 & add126_376 & add135_401;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1119_inst WPIPE_Block3_start_1122_inst WPIPE_Block3_start_1125_inst WPIPE_Block3_start_1128_inst WPIPE_Block3_start_1131_inst WPIPE_Block3_start_1134_inst WPIPE_Block3_start_1137_inst WPIPE_Block3_start_1140_inst WPIPE_Block3_start_1143_inst WPIPE_Block3_start_1156_inst WPIPE_Block3_start_1163_inst WPIPE_Block3_start_1166_inst WPIPE_Block3_start_1169_inst WPIPE_Block3_start_1172_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1119_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1122_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1125_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1128_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1131_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1134_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1137_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1140_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1143_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1156_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1163_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1166_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1169_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1172_inst_req_0;
      WPIPE_Block3_start_1119_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1122_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1125_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1128_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1131_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1134_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1137_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1140_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1143_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1156_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1163_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1166_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1169_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1172_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1119_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1122_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1125_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1128_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1131_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1134_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1137_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1140_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1143_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1156_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1163_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1166_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1169_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1172_inst_req_1;
      WPIPE_Block3_start_1119_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1122_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1125_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1128_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1131_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1134_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1137_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1140_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1143_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1156_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1163_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1166_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1169_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1172_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_50 & add12_75 & add21_100 & add30_125 & add39_150 & add48_175 & add57_200 & add99_301 & add108_326 & conv336_1155 & conv338_1162 & add117_351 & add126_376 & add135_401;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1355_inst WPIPE_ConvTranspose_output_pipe_1349_inst WPIPE_ConvTranspose_output_pipe_1352_inst WPIPE_ConvTranspose_output_pipe_1334_inst WPIPE_ConvTranspose_output_pipe_1337_inst WPIPE_ConvTranspose_output_pipe_1340_inst WPIPE_ConvTranspose_output_pipe_1343_inst WPIPE_ConvTranspose_output_pipe_1346_inst WPIPE_ConvTranspose_output_pipe_954_inst WPIPE_ConvTranspose_output_pipe_958_inst WPIPE_ConvTranspose_output_pipe_1188_inst WPIPE_ConvTranspose_output_pipe_1192_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1355_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1349_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1352_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1334_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1337_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1340_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1343_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1346_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_954_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_958_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1188_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1192_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1355_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1349_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1352_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1334_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1337_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1340_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1343_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1346_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_954_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_958_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1188_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1192_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1355_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1349_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1352_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1334_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1337_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1340_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1343_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1346_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_954_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_958_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1188_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1192_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1355_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1349_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1352_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1334_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1337_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1340_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1343_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1346_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_954_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_958_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1188_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1192_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= conv365_1263 & conv377_1283 & conv371_1273 & conv407_1333 & conv401_1323 & conv395_1313 & conv389_1303 & conv383_1293 & type_cast_956_wire_constant & type_cast_960_wire_constant & type_cast_1190_wire_constant & type_cast_1194_wire_constant;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3500_start: Boolean;
  signal convTransposeA_CP_3500_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_start_1443_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1425_inst_ack_1 : boolean;
  signal array_obj_ref_1598_index_offset_ack_1 : boolean;
  signal array_obj_ref_1598_index_offset_req_1 : boolean;
  signal type_cast_1482_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1437_inst_ack_1 : boolean;
  signal type_cast_1592_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1440_inst_req_0 : boolean;
  signal type_cast_1592_inst_ack_0 : boolean;
  signal type_cast_1630_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1437_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1443_inst_req_1 : boolean;
  signal addr_of_1599_final_reg_req_1 : boolean;
  signal ptr_deref_1625_store_0_ack_1 : boolean;
  signal RPIPE_Block0_start_1425_inst_req_1 : boolean;
  signal addr_of_1622_final_reg_ack_0 : boolean;
  signal type_cast_1482_inst_req_0 : boolean;
  signal type_cast_1592_inst_req_0 : boolean;
  signal type_cast_1482_inst_ack_0 : boolean;
  signal array_obj_ref_1621_index_offset_req_1 : boolean;
  signal addr_of_1622_final_reg_req_0 : boolean;
  signal type_cast_1482_inst_ack_1 : boolean;
  signal type_cast_1630_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1437_inst_ack_0 : boolean;
  signal array_obj_ref_1621_index_offset_ack_1 : boolean;
  signal array_obj_ref_1621_index_offset_ack_0 : boolean;
  signal type_cast_1478_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1425_inst_ack_0 : boolean;
  signal ptr_deref_1625_store_0_ack_0 : boolean;
  signal RPIPE_Block0_start_1425_inst_req_0 : boolean;
  signal type_cast_1478_inst_req_1 : boolean;
  signal array_obj_ref_1598_index_offset_ack_0 : boolean;
  signal array_obj_ref_1598_index_offset_req_0 : boolean;
  signal type_cast_1478_inst_ack_0 : boolean;
  signal type_cast_1478_inst_req_0 : boolean;
  signal addr_of_1599_final_reg_ack_1 : boolean;
  signal RPIPE_Block0_start_1440_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1437_inst_req_0 : boolean;
  signal array_obj_ref_1621_index_offset_req_0 : boolean;
  signal type_cast_1554_inst_req_1 : boolean;
  signal type_cast_1630_inst_ack_1 : boolean;
  signal addr_of_1599_final_reg_req_0 : boolean;
  signal type_cast_1558_inst_ack_1 : boolean;
  signal addr_of_1622_final_reg_req_1 : boolean;
  signal addr_of_1599_final_reg_ack_0 : boolean;
  signal type_cast_1558_inst_req_0 : boolean;
  signal type_cast_1592_inst_ack_1 : boolean;
  signal ptr_deref_1625_store_0_req_0 : boolean;
  signal addr_of_1622_final_reg_ack_1 : boolean;
  signal if_stmt_1643_branch_ack_0 : boolean;
  signal ptr_deref_1603_load_0_ack_1 : boolean;
  signal type_cast_1416_inst_ack_1 : boolean;
  signal ptr_deref_1603_load_0_req_1 : boolean;
  signal if_stmt_1643_branch_req_0 : boolean;
  signal type_cast_1554_inst_ack_0 : boolean;
  signal type_cast_1671_inst_req_0 : boolean;
  signal type_cast_1671_inst_ack_0 : boolean;
  signal type_cast_1554_inst_req_0 : boolean;
  signal type_cast_1671_inst_ack_1 : boolean;
  signal type_cast_1554_inst_ack_1 : boolean;
  signal ptr_deref_1603_load_0_req_0 : boolean;
  signal type_cast_1671_inst_req_1 : boolean;
  signal if_stmt_1643_branch_ack_1 : boolean;
  signal ptr_deref_1603_load_0_ack_0 : boolean;
  signal type_cast_1558_inst_ack_0 : boolean;
  signal type_cast_1470_inst_req_0 : boolean;
  signal type_cast_1630_inst_ack_0 : boolean;
  signal ptr_deref_1625_store_0_req_1 : boolean;
  signal type_cast_1558_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1443_inst_ack_0 : boolean;
  signal type_cast_1470_inst_ack_1 : boolean;
  signal type_cast_1416_inst_req_1 : boolean;
  signal type_cast_1470_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1443_inst_req_0 : boolean;
  signal type_cast_1470_inst_ack_0 : boolean;
  signal type_cast_1562_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1385_inst_req_0 : boolean;
  signal type_cast_1562_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1385_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1385_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1385_inst_ack_1 : boolean;
  signal type_cast_1474_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1388_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1388_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1388_inst_req_1 : boolean;
  signal type_cast_1562_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1388_inst_ack_1 : boolean;
  signal type_cast_1474_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1391_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1391_inst_ack_0 : boolean;
  signal type_cast_1562_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1391_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1391_inst_ack_1 : boolean;
  signal type_cast_1429_inst_ack_1 : boolean;
  signal type_cast_1429_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1394_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1394_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1394_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1394_inst_ack_1 : boolean;
  signal type_cast_1429_inst_ack_0 : boolean;
  signal type_cast_1429_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1397_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1397_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1440_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1397_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1397_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1440_inst_req_1 : boolean;
  signal type_cast_1474_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1400_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1400_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1400_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1400_inst_ack_1 : boolean;
  signal type_cast_1474_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1403_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1403_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1403_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1403_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1406_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1406_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1406_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1406_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1409_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1409_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1409_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1409_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1412_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1412_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1412_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1412_inst_ack_1 : boolean;
  signal type_cast_1416_inst_req_0 : boolean;
  signal type_cast_1416_inst_ack_0 : boolean;
  signal type_cast_1687_inst_req_0 : boolean;
  signal type_cast_1687_inst_ack_0 : boolean;
  signal type_cast_1687_inst_req_1 : boolean;
  signal type_cast_1687_inst_ack_1 : boolean;
  signal if_stmt_1694_branch_req_0 : boolean;
  signal if_stmt_1694_branch_ack_1 : boolean;
  signal if_stmt_1694_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1730_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1730_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1730_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1730_inst_ack_1 : boolean;
  signal phi_stmt_1492_req_0 : boolean;
  signal phi_stmt_1499_req_0 : boolean;
  signal phi_stmt_1506_req_0 : boolean;
  signal phi_stmt_1513_req_0 : boolean;
  signal type_cast_1498_inst_req_0 : boolean;
  signal type_cast_1498_inst_ack_0 : boolean;
  signal type_cast_1498_inst_req_1 : boolean;
  signal type_cast_1498_inst_ack_1 : boolean;
  signal phi_stmt_1492_req_1 : boolean;
  signal type_cast_1505_inst_req_0 : boolean;
  signal type_cast_1505_inst_ack_0 : boolean;
  signal type_cast_1505_inst_req_1 : boolean;
  signal type_cast_1505_inst_ack_1 : boolean;
  signal phi_stmt_1499_req_1 : boolean;
  signal type_cast_1512_inst_req_0 : boolean;
  signal type_cast_1512_inst_ack_0 : boolean;
  signal type_cast_1512_inst_req_1 : boolean;
  signal type_cast_1512_inst_ack_1 : boolean;
  signal phi_stmt_1506_req_1 : boolean;
  signal type_cast_1519_inst_req_0 : boolean;
  signal type_cast_1519_inst_ack_0 : boolean;
  signal type_cast_1519_inst_req_1 : boolean;
  signal type_cast_1519_inst_ack_1 : boolean;
  signal phi_stmt_1513_req_1 : boolean;
  signal phi_stmt_1492_ack_0 : boolean;
  signal phi_stmt_1499_ack_0 : boolean;
  signal phi_stmt_1506_ack_0 : boolean;
  signal phi_stmt_1513_ack_0 : boolean;
  signal phi_stmt_1701_req_1 : boolean;
  signal type_cast_1713_inst_req_0 : boolean;
  signal type_cast_1713_inst_ack_0 : boolean;
  signal type_cast_1713_inst_req_1 : boolean;
  signal type_cast_1713_inst_ack_1 : boolean;
  signal phi_stmt_1708_req_1 : boolean;
  signal type_cast_1719_inst_req_0 : boolean;
  signal type_cast_1719_inst_ack_0 : boolean;
  signal type_cast_1719_inst_req_1 : boolean;
  signal type_cast_1719_inst_ack_1 : boolean;
  signal phi_stmt_1714_req_1 : boolean;
  signal type_cast_1704_inst_req_0 : boolean;
  signal type_cast_1704_inst_ack_0 : boolean;
  signal type_cast_1704_inst_req_1 : boolean;
  signal type_cast_1704_inst_ack_1 : boolean;
  signal phi_stmt_1701_req_0 : boolean;
  signal type_cast_1711_inst_req_0 : boolean;
  signal type_cast_1711_inst_ack_0 : boolean;
  signal type_cast_1711_inst_req_1 : boolean;
  signal type_cast_1711_inst_ack_1 : boolean;
  signal phi_stmt_1708_req_0 : boolean;
  signal type_cast_1717_inst_req_0 : boolean;
  signal type_cast_1717_inst_ack_0 : boolean;
  signal type_cast_1717_inst_req_1 : boolean;
  signal type_cast_1717_inst_ack_1 : boolean;
  signal phi_stmt_1714_req_0 : boolean;
  signal phi_stmt_1701_ack_0 : boolean;
  signal phi_stmt_1708_ack_0 : boolean;
  signal phi_stmt_1714_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3500_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3500_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3500_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3500_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3500: Block -- control-path 
    signal convTransposeA_CP_3500_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3500_elements(0) <= convTransposeA_CP_3500_start;
    convTransposeA_CP_3500_symbol <= convTransposeA_CP_3500_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1383/$entry
      -- CP-element group 0: 	 branch_block_stmt_1383/branch_block_stmt_1383__entry__
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444__entry__
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/$entry
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_update_start_
      -- 
    cr_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(0), ack => type_cast_1416_inst_req_1); -- 
    rr_3548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(0), ack => RPIPE_Block0_start_1385_inst_req_0); -- 
    cr_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(0), ack => type_cast_1429_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1383/merge_stmt_1700__exit__
      -- CP-element group 1: 	 branch_block_stmt_1383/assign_stmt_1726__entry__
      -- CP-element group 1: 	 branch_block_stmt_1383/assign_stmt_1726__exit__
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1383/assign_stmt_1726/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/assign_stmt_1726/$exit
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/cr
      -- 
    rr_4234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1498_inst_req_0); -- 
    cr_4239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1498_inst_req_1); -- 
    rr_4257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1505_inst_req_0); -- 
    cr_4262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1505_inst_req_1); -- 
    rr_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1512_inst_req_0); -- 
    cr_4285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1512_inst_req_1); -- 
    rr_4303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1519_inst_req_0); -- 
    cr_4308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(1), ack => type_cast_1519_inst_req_1); -- 
    convTransposeA_CP_3500_elements(1) <= convTransposeA_CP_3500_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Update/cr
      -- 
    ra_3549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1385_inst_ack_0, ack => convTransposeA_CP_3500_elements(2)); -- 
    cr_3553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(2), ack => RPIPE_Block0_start_1385_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1385_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Sample/rr
      -- 
    ca_3554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1385_inst_ack_1, ack => convTransposeA_CP_3500_elements(3)); -- 
    rr_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(3), ack => RPIPE_Block0_start_1388_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Update/cr
      -- 
    ra_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1388_inst_ack_0, ack => convTransposeA_CP_3500_elements(4)); -- 
    cr_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(4), ack => RPIPE_Block0_start_1388_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1388_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Sample/rr
      -- 
    ca_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1388_inst_ack_1, ack => convTransposeA_CP_3500_elements(5)); -- 
    rr_3576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(5), ack => RPIPE_Block0_start_1391_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Update/cr
      -- 
    ra_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1391_inst_ack_0, ack => convTransposeA_CP_3500_elements(6)); -- 
    cr_3581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(6), ack => RPIPE_Block0_start_1391_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1391_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Sample/rr
      -- 
    ca_3582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1391_inst_ack_1, ack => convTransposeA_CP_3500_elements(7)); -- 
    rr_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(7), ack => RPIPE_Block0_start_1394_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Update/cr
      -- 
    ra_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1394_inst_ack_0, ack => convTransposeA_CP_3500_elements(8)); -- 
    cr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(8), ack => RPIPE_Block0_start_1394_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1394_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Sample/rr
      -- 
    ca_3596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1394_inst_ack_1, ack => convTransposeA_CP_3500_elements(9)); -- 
    rr_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(9), ack => RPIPE_Block0_start_1397_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Update/cr
      -- 
    ra_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1397_inst_ack_0, ack => convTransposeA_CP_3500_elements(10)); -- 
    cr_3609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(10), ack => RPIPE_Block0_start_1397_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1397_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Sample/rr
      -- 
    ca_3610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1397_inst_ack_1, ack => convTransposeA_CP_3500_elements(11)); -- 
    rr_3618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(11), ack => RPIPE_Block0_start_1400_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Update/cr
      -- 
    ra_3619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1400_inst_ack_0, ack => convTransposeA_CP_3500_elements(12)); -- 
    cr_3623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(12), ack => RPIPE_Block0_start_1400_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1400_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Sample/rr
      -- 
    ca_3624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1400_inst_ack_1, ack => convTransposeA_CP_3500_elements(13)); -- 
    rr_3632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(13), ack => RPIPE_Block0_start_1403_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Update/cr
      -- 
    ra_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1403_inst_ack_0, ack => convTransposeA_CP_3500_elements(14)); -- 
    cr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(14), ack => RPIPE_Block0_start_1403_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1403_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Sample/rr
      -- 
    ca_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1403_inst_ack_1, ack => convTransposeA_CP_3500_elements(15)); -- 
    rr_3646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(15), ack => RPIPE_Block0_start_1406_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Update/cr
      -- 
    ra_3647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1406_inst_ack_0, ack => convTransposeA_CP_3500_elements(16)); -- 
    cr_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(16), ack => RPIPE_Block0_start_1406_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1406_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Sample/rr
      -- 
    ca_3652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1406_inst_ack_1, ack => convTransposeA_CP_3500_elements(17)); -- 
    rr_3660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(17), ack => RPIPE_Block0_start_1409_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Update/cr
      -- 
    ra_3661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1409_inst_ack_0, ack => convTransposeA_CP_3500_elements(18)); -- 
    cr_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(18), ack => RPIPE_Block0_start_1409_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1409_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Sample/rr
      -- 
    ca_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1409_inst_ack_1, ack => convTransposeA_CP_3500_elements(19)); -- 
    rr_3674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(19), ack => RPIPE_Block0_start_1412_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Update/cr
      -- 
    ra_3675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1412_inst_ack_0, ack => convTransposeA_CP_3500_elements(20)); -- 
    cr_3679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(20), ack => RPIPE_Block0_start_1412_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1412_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Sample/rr
      -- 
    ca_3680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1412_inst_ack_1, ack => convTransposeA_CP_3500_elements(21)); -- 
    rr_3688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(21), ack => type_cast_1416_inst_req_0); -- 
    rr_3702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(21), ack => RPIPE_Block0_start_1425_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Sample/ra
      -- 
    ra_3689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_0, ack => convTransposeA_CP_3500_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1416_update_completed_
      -- 
    ca_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_1, ack => convTransposeA_CP_3500_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_sample_completed_
      -- 
    ra_3703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1425_inst_ack_0, ack => convTransposeA_CP_3500_elements(24)); -- 
    cr_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(24), ack => RPIPE_Block0_start_1425_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1425_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Sample/$entry
      -- 
    ca_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1425_inst_ack_1, ack => convTransposeA_CP_3500_elements(25)); -- 
    rr_3716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(25), ack => type_cast_1429_inst_req_0); -- 
    rr_3730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(25), ack => RPIPE_Block0_start_1437_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Sample/$exit
      -- 
    ra_3717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_0, ack => convTransposeA_CP_3500_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/type_cast_1429_update_completed_
      -- 
    ca_3722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_1, ack => convTransposeA_CP_3500_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_sample_completed_
      -- 
    ra_3731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1437_inst_ack_0, ack => convTransposeA_CP_3500_elements(28)); -- 
    cr_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(28), ack => RPIPE_Block0_start_1437_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1437_update_completed_
      -- 
    ca_3736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1437_inst_ack_1, ack => convTransposeA_CP_3500_elements(29)); -- 
    rr_3744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(29), ack => RPIPE_Block0_start_1440_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Update/$entry
      -- 
    ra_3745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1440_inst_ack_0, ack => convTransposeA_CP_3500_elements(30)); -- 
    cr_3749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(30), ack => RPIPE_Block0_start_1440_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1440_Update/$exit
      -- 
    ca_3750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1440_inst_ack_1, ack => convTransposeA_CP_3500_elements(31)); -- 
    rr_3758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(31), ack => RPIPE_Block0_start_1443_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_sample_completed_
      -- 
    ra_3759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1443_inst_ack_0, ack => convTransposeA_CP_3500_elements(32)); -- 
    cr_3763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(32), ack => RPIPE_Block0_start_1443_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/RPIPE_Block0_start_1443_update_completed_
      -- 
    ca_3764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1443_inst_ack_1, ack => convTransposeA_CP_3500_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444__exit__
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489__entry__
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1386_to_assign_stmt_1444/$exit
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Sample/rr
      -- 
    cr_3822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1482_inst_req_1); -- 
    rr_3817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1482_inst_req_0); -- 
    cr_3808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1478_inst_req_1); -- 
    rr_3803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1478_inst_req_0); -- 
    rr_3775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1470_inst_req_0); -- 
    cr_3780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1470_inst_req_1); -- 
    cr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1474_inst_req_1); -- 
    rr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(34), ack => type_cast_1474_inst_req_0); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(23) & convTransposeA_CP_3500_elements(27) & convTransposeA_CP_3500_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Sample/ra
      -- 
    ra_3776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1470_inst_ack_0, ack => convTransposeA_CP_3500_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1470_Update/$exit
      -- 
    ca_3781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1470_inst_ack_1, ack => convTransposeA_CP_3500_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Sample/ra
      -- 
    ra_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1474_inst_ack_0, ack => convTransposeA_CP_3500_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1474_Update/$exit
      -- 
    ca_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1474_inst_ack_1, ack => convTransposeA_CP_3500_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Sample/$exit
      -- 
    ra_3804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1478_inst_ack_0, ack => convTransposeA_CP_3500_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1478_Update/$exit
      -- 
    ca_3809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1478_inst_ack_1, ack => convTransposeA_CP_3500_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_sample_completed_
      -- 
    ra_3818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1482_inst_ack_0, ack => convTransposeA_CP_3500_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/type_cast_1482_Update/ca
      -- 
    ca_3823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1482_inst_ack_1, ack => convTransposeA_CP_3500_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489/$exit
      -- CP-element group 43: 	 branch_block_stmt_1383/assign_stmt_1451_to_assign_stmt_1489__exit__
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1492/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1499/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1506/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1513/$entry
      -- CP-element group 43: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(36) & convTransposeA_CP_3500_elements(38) & convTransposeA_CP_3500_elements(40) & convTransposeA_CP_3500_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_sample_completed_
      -- 
    ra_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_0, ack => convTransposeA_CP_3500_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Update/ca
      -- 
    ca_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_1, ack => convTransposeA_CP_3500_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Sample/ra
      -- 
    ra_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1558_inst_ack_0, ack => convTransposeA_CP_3500_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Update/$exit
      -- 
    ca_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1558_inst_ack_1, ack => convTransposeA_CP_3500_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_sample_completed_
      -- 
    ra_3863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1562_inst_ack_0, ack => convTransposeA_CP_3500_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_update_completed_
      -- 
    ca_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1562_inst_ack_1, ack => convTransposeA_CP_3500_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_sample_completed_
      -- 
    ra_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_0, ack => convTransposeA_CP_3500_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_index_resize_1/index_resize_ack
      -- 
    ca_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_1, ack => convTransposeA_CP_3500_elements(51)); -- 
    req_3907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(51), ack => array_obj_ref_1598_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Sample/$exit
      -- 
    ack_3908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1598_index_offset_ack_0, ack => convTransposeA_CP_3500_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_request/req
      -- CP-element group 53: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_request/$entry
      -- 
    ack_3913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1598_index_offset_ack_1, ack => convTransposeA_CP_3500_elements(53)); -- 
    req_3922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(53), ack => addr_of_1599_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_request/ack
      -- CP-element group 54: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_request/$exit
      -- 
    ack_3923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1599_final_reg_ack_0, ack => convTransposeA_CP_3500_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/word_access_start/word_0/rr
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_base_address_resized
      -- 
    ack_3928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1599_final_reg_ack_1, ack => convTransposeA_CP_3500_elements(55)); -- 
    rr_3961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(55), ack => ptr_deref_1603_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Sample/word_access_start/word_0/ra
      -- 
    ra_3962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1603_load_0_ack_0, ack => convTransposeA_CP_3500_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/ptr_deref_1603_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/ptr_deref_1603_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/ptr_deref_1603_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/ptr_deref_1603_Merge/merge_ack
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/word_access_complete/$exit
      -- 
    ca_3973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1603_load_0_ack_1, ack => convTransposeA_CP_3500_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_index_resized_1
      -- 
    req_4003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(58), ack => array_obj_ref_1621_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(45) & convTransposeA_CP_3500_elements(47) & convTransposeA_CP_3500_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_sample_complete
      -- 
    ack_4004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1621_index_offset_ack_0, ack => convTransposeA_CP_3500_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_request/req
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_root_address_calculated
      -- 
    ack_4009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1621_index_offset_ack_1, ack => convTransposeA_CP_3500_elements(60)); -- 
    req_4018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(60), ack => addr_of_1622_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_request/ack
      -- 
    ack_4019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1622_final_reg_ack_0, ack => convTransposeA_CP_3500_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_update_completed_
      -- 
    ack_4024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1622_final_reg_ack_1, ack => convTransposeA_CP_3500_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/ptr_deref_1625_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/ptr_deref_1625_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/ptr_deref_1625_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/ptr_deref_1625_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/word_access_start/word_0/rr
      -- CP-element group 63: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_sample_start_
      -- 
    rr_4062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(63), ack => ptr_deref_1625_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(57) & convTransposeA_CP_3500_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/word_access_start/word_0/ra
      -- CP-element group 64: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_sample_completed_
      -- 
    ra_4063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1625_store_0_ack_0, ack => convTransposeA_CP_3500_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/word_access_complete/word_0/ca
      -- CP-element group 65: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_update_completed_
      -- 
    ca_4074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1625_store_0_ack_1, ack => convTransposeA_CP_3500_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Sample/ra
      -- 
    ra_4083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1630_inst_ack_0, ack => convTransposeA_CP_3500_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Update/$exit
      -- 
    ca_4088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1630_inst_ack_1, ack => convTransposeA_CP_3500_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/$exit
      -- CP-element group 68: 	 branch_block_stmt_1383/if_stmt_1643_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1383/if_stmt_1643_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1383/if_stmt_1643_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1383/if_stmt_1643_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1383/if_stmt_1643_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1383/if_stmt_1643_else_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642__exit__
      -- CP-element group 68: 	 branch_block_stmt_1383/if_stmt_1643__entry__
      -- CP-element group 68: 	 branch_block_stmt_1383/R_cmp_1644_place
      -- 
    branch_req_4096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(68), ack => if_stmt_1643_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(52) & convTransposeA_CP_3500_elements(59) & convTransposeA_CP_3500_elements(65) & convTransposeA_CP_3500_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1383/assign_stmt_1655/$exit
      -- CP-element group 69: 	 branch_block_stmt_1383/if_stmt_1643_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1383/if_stmt_1643_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1383/assign_stmt_1655/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/merge_stmt_1649__exit__
      -- CP-element group 69: 	 branch_block_stmt_1383/assign_stmt_1655__entry__
      -- CP-element group 69: 	 branch_block_stmt_1383/assign_stmt_1655__exit__
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1383/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1383/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1383/merge_stmt_1649_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1383/merge_stmt_1649_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/merge_stmt_1649_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1383/merge_stmt_1649_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1643_branch_ack_1, ack => convTransposeA_CP_3500_elements(69)); -- 
    rr_4418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(69), ack => type_cast_1704_inst_req_0); -- 
    cr_4423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(69), ack => type_cast_1704_inst_req_1); -- 
    rr_4441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(69), ack => type_cast_1711_inst_req_0); -- 
    cr_4446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(69), ack => type_cast_1711_inst_req_1); -- 
    rr_4464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(69), ack => type_cast_1717_inst_req_0); -- 
    cr_4469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(69), ack => type_cast_1717_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1383/if_stmt_1643_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/$entry
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1383/if_stmt_1643_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1383/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1383/merge_stmt_1657__exit__
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693__entry__
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1383/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1383/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1383/merge_stmt_1657_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1383/merge_stmt_1657_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1383/merge_stmt_1657_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1383/merge_stmt_1657_PhiAck/dummy
      -- 
    else_choice_transition_4105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1643_branch_ack_0, ack => convTransposeA_CP_3500_elements(70)); -- 
    rr_4121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(70), ack => type_cast_1671_inst_req_0); -- 
    cr_4126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(70), ack => type_cast_1671_inst_req_1); -- 
    cr_4140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(70), ack => type_cast_1687_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Sample/ra
      -- 
    ra_4122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_0, ack => convTransposeA_CP_3500_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1671_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Sample/rr
      -- 
    ca_4127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_1, ack => convTransposeA_CP_3500_elements(72)); -- 
    rr_4135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(72), ack => type_cast_1687_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Sample/ra
      -- 
    ra_4136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1687_inst_ack_0, ack => convTransposeA_CP_3500_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/$exit
      -- CP-element group 74: 	 branch_block_stmt_1383/R_cmp112_1695_place
      -- CP-element group 74: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693__exit__
      -- CP-element group 74: 	 branch_block_stmt_1383/if_stmt_1694__entry__
      -- CP-element group 74: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1383/assign_stmt_1663_to_assign_stmt_1693/type_cast_1687_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1383/if_stmt_1694_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1383/if_stmt_1694_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1383/if_stmt_1694_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1383/if_stmt_1694_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1383/if_stmt_1694_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1383/if_stmt_1694_else_link/$entry
      -- 
    ca_4141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1687_inst_ack_1, ack => convTransposeA_CP_3500_elements(74)); -- 
    branch_req_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(74), ack => if_stmt_1694_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1383/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1383/merge_stmt_1728__exit__
      -- CP-element group 75: 	 branch_block_stmt_1383/assign_stmt_1733__entry__
      -- CP-element group 75: 	 branch_block_stmt_1383/if_stmt_1694_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1383/if_stmt_1694_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1383/assign_stmt_1733/$entry
      -- CP-element group 75: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1383/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1383/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1383/merge_stmt_1728_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1383/merge_stmt_1728_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1383/merge_stmt_1728_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1383/merge_stmt_1728_PhiAck/dummy
      -- 
    if_choice_transition_4154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1694_branch_ack_1, ack => convTransposeA_CP_3500_elements(75)); -- 
    req_4174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(75), ack => WPIPE_Block0_done_1730_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	108 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123
      -- CP-element group 76: 	 branch_block_stmt_1383/if_stmt_1694_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1383/if_stmt_1694_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1701/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1694_branch_ack_0, ack => convTransposeA_CP_3500_elements(76)); -- 
    rr_4369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(76), ack => type_cast_1713_inst_req_0); -- 
    cr_4374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(76), ack => type_cast_1713_inst_req_1); -- 
    rr_4392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(76), ack => type_cast_1719_inst_req_0); -- 
    cr_4397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(76), ack => type_cast_1719_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Update/req
      -- 
    ack_4175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1730_inst_ack_0, ack => convTransposeA_CP_3500_elements(77)); -- 
    req_4179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(77), ack => WPIPE_Block0_done_1730_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1383/$exit
      -- CP-element group 78: 	 branch_block_stmt_1383/branch_block_stmt_1383__exit__
      -- CP-element group 78: 	 branch_block_stmt_1383/assign_stmt_1733__exit__
      -- CP-element group 78: 	 branch_block_stmt_1383/return__
      -- CP-element group 78: 	 branch_block_stmt_1383/merge_stmt_1735__exit__
      -- CP-element group 78: 	 branch_block_stmt_1383/assign_stmt_1733/$exit
      -- CP-element group 78: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1383/assign_stmt_1733/WPIPE_Block0_done_1730_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1383/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1383/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1383/merge_stmt_1735_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1383/merge_stmt_1735_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1383/merge_stmt_1735_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1383/merge_stmt_1735_PhiAck/dummy
      -- 
    ack_4180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1730_inst_ack_1, ack => convTransposeA_CP_3500_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1492/$exit
      -- CP-element group 79: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1496_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_req
      -- 
    phi_stmt_1492_req_4191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1492_req_4191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(79), ack => phi_stmt_1492_req_0); -- 
    -- Element group convTransposeA_CP_3500_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3500_elements(43), ack => convTransposeA_CP_3500_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1499/$exit
      -- CP-element group 80: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1503_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_req
      -- 
    phi_stmt_1499_req_4199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1499_req_4199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(80), ack => phi_stmt_1499_req_0); -- 
    -- Element group convTransposeA_CP_3500_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3500_elements(43), ack => convTransposeA_CP_3500_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1506/$exit
      -- CP-element group 81: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1510_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_req
      -- 
    phi_stmt_1506_req_4207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1506_req_4207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(81), ack => phi_stmt_1506_req_0); -- 
    -- Element group convTransposeA_CP_3500_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3500_elements(43), ack => convTransposeA_CP_3500_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1513/$exit
      -- CP-element group 82: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1517_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_req
      -- 
    phi_stmt_1513_req_4215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1513_req_4215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(82), ack => phi_stmt_1513_req_0); -- 
    -- Element group convTransposeA_CP_3500_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3500_elements(43), ack => convTransposeA_CP_3500_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1383/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(79) & convTransposeA_CP_3500_elements(80) & convTransposeA_CP_3500_elements(81) & convTransposeA_CP_3500_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Sample/ra
      -- 
    ra_4235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1498_inst_ack_0, ack => convTransposeA_CP_3500_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/Update/ca
      -- 
    ca_4240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1498_inst_ack_1, ack => convTransposeA_CP_3500_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/$exit
      -- CP-element group 86: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/$exit
      -- CP-element group 86: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_sources/type_cast_1498/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1492/phi_stmt_1492_req
      -- 
    phi_stmt_1492_req_4241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1492_req_4241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(86), ack => phi_stmt_1492_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(84) & convTransposeA_CP_3500_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Sample/ra
      -- 
    ra_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1505_inst_ack_0, ack => convTransposeA_CP_3500_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/Update/ca
      -- 
    ca_4263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1505_inst_ack_1, ack => convTransposeA_CP_3500_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/$exit
      -- CP-element group 89: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/$exit
      -- CP-element group 89: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_sources/type_cast_1505/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1499/phi_stmt_1499_req
      -- 
    phi_stmt_1499_req_4264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1499_req_4264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(89), ack => phi_stmt_1499_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(87) & convTransposeA_CP_3500_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/ra
      -- 
    ra_4281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1512_inst_ack_0, ack => convTransposeA_CP_3500_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/ca
      -- 
    ca_4286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1512_inst_ack_1, ack => convTransposeA_CP_3500_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/$exit
      -- CP-element group 92: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/$exit
      -- CP-element group 92: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_req
      -- 
    phi_stmt_1506_req_4287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1506_req_4287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(92), ack => phi_stmt_1506_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(90) & convTransposeA_CP_3500_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/ra
      -- 
    ra_4304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1519_inst_ack_0, ack => convTransposeA_CP_3500_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/ca
      -- 
    ca_4309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1519_inst_ack_1, ack => convTransposeA_CP_3500_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/$exit
      -- CP-element group 95: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/$exit
      -- CP-element group 95: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_req
      -- 
    phi_stmt_1513_req_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1513_req_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(95), ack => phi_stmt_1513_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(93) & convTransposeA_CP_3500_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1383/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(86) & convTransposeA_CP_3500_elements(89) & convTransposeA_CP_3500_elements(92) & convTransposeA_CP_3500_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1383/merge_stmt_1491_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_1383/merge_stmt_1491_PhiAck/$entry
      -- 
    convTransposeA_CP_3500_elements(97) <= OrReduce(convTransposeA_CP_3500_elements(83) & convTransposeA_CP_3500_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1383/merge_stmt_1491_PhiAck/phi_stmt_1492_ack
      -- 
    phi_stmt_1492_ack_4315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1492_ack_0, ack => convTransposeA_CP_3500_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1383/merge_stmt_1491_PhiAck/phi_stmt_1499_ack
      -- 
    phi_stmt_1499_ack_4316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1499_ack_0, ack => convTransposeA_CP_3500_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1383/merge_stmt_1491_PhiAck/phi_stmt_1506_ack
      -- 
    phi_stmt_1506_ack_4317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1506_ack_0, ack => convTransposeA_CP_3500_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1383/merge_stmt_1491_PhiAck/phi_stmt_1513_ack
      -- 
    phi_stmt_1513_ack_4318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1513_ack_0, ack => convTransposeA_CP_3500_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1599_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1598_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1630_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1554_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1603_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/ptr_deref_1625_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1558_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1592_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/merge_stmt_1491__exit__
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642__entry__
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/array_obj_ref_1621_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/type_cast_1562_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/assign_stmt_1526_to_assign_stmt_1642/addr_of_1622_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1383/merge_stmt_1491_PhiAck/$exit
      -- 
    req_3912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => array_obj_ref_1598_index_offset_req_1); -- 
    cr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1592_inst_req_1); -- 
    cr_4087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1630_inst_req_1); -- 
    req_3927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => addr_of_1599_final_reg_req_1); -- 
    rr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1592_inst_req_0); -- 
    req_4008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => array_obj_ref_1621_index_offset_req_1); -- 
    rr_4082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1630_inst_req_0); -- 
    cr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1554_inst_req_1); -- 
    req_4023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => addr_of_1622_final_reg_req_1); -- 
    rr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1558_inst_req_0); -- 
    cr_3972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => ptr_deref_1603_load_0_req_1); -- 
    rr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1554_inst_req_0); -- 
    cr_4073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => ptr_deref_1625_store_0_req_1); -- 
    cr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1558_inst_req_1); -- 
    cr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1562_inst_req_1); -- 
    rr_3862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(102), ack => type_cast_1562_inst_req_0); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(98) & convTransposeA_CP_3500_elements(99) & convTransposeA_CP_3500_elements(100) & convTransposeA_CP_3500_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  output  delay-element  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	110 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1701/$exit
      -- CP-element group 103: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1707_konst_delay_trans
      -- CP-element group 103: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_req
      -- 
    phi_stmt_1701_req_4353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1701_req_4353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(103), ack => phi_stmt_1701_req_1); -- 
    -- Element group convTransposeA_CP_3500_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => convTransposeA_CP_3500_elements(76), ack => convTransposeA_CP_3500_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Sample/ra
      -- 
    ra_4370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1713_inst_ack_0, ack => convTransposeA_CP_3500_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/Update/ca
      -- 
    ca_4375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1713_inst_ack_1, ack => convTransposeA_CP_3500_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/$exit
      -- CP-element group 106: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/$exit
      -- CP-element group 106: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/$exit
      -- CP-element group 106: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1713/SplitProtocol/$exit
      -- CP-element group 106: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_req
      -- 
    phi_stmt_1708_req_4376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1708_req_4376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(106), ack => phi_stmt_1708_req_1); -- 
    convTransposeA_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(104) & convTransposeA_CP_3500_elements(105);
      gj_convTransposeA_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Sample/ra
      -- 
    ra_4393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1719_inst_ack_0, ack => convTransposeA_CP_3500_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/Update/ca
      -- 
    ca_4398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1719_inst_ack_1, ack => convTransposeA_CP_3500_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/$exit
      -- CP-element group 109: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/$exit
      -- CP-element group 109: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1719/SplitProtocol/$exit
      -- CP-element group 109: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_req
      -- 
    phi_stmt_1714_req_4399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1714_req_4399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(109), ack => phi_stmt_1714_req_1); -- 
    convTransposeA_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(107) & convTransposeA_CP_3500_elements(108);
      gj_convTransposeA_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1383/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(103) & convTransposeA_CP_3500_elements(106) & convTransposeA_CP_3500_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Sample/ra
      -- 
    ra_4419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1704_inst_ack_0, ack => convTransposeA_CP_3500_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/Update/ca
      -- 
    ca_4424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1704_inst_ack_1, ack => convTransposeA_CP_3500_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/$exit
      -- CP-element group 113: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/$exit
      -- CP-element group 113: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_sources/type_cast_1704/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1701/phi_stmt_1701_req
      -- 
    phi_stmt_1701_req_4425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1701_req_4425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(113), ack => phi_stmt_1701_req_0); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(111) & convTransposeA_CP_3500_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Sample/ra
      -- 
    ra_4442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_0, ack => convTransposeA_CP_3500_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/Update/ca
      -- 
    ca_4447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_1, ack => convTransposeA_CP_3500_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/$exit
      -- CP-element group 116: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/$exit
      -- CP-element group 116: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_sources/type_cast_1711/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1708/phi_stmt_1708_req
      -- 
    phi_stmt_1708_req_4448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1708_req_4448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(116), ack => phi_stmt_1708_req_0); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(114) & convTransposeA_CP_3500_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Sample/ra
      -- 
    ra_4465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1717_inst_ack_0, ack => convTransposeA_CP_3500_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/Update/ca
      -- 
    ca_4470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1717_inst_ack_1, ack => convTransposeA_CP_3500_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/$exit
      -- CP-element group 119: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/$exit
      -- CP-element group 119: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_sources/type_cast_1717/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1714/phi_stmt_1714_req
      -- 
    phi_stmt_1714_req_4471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1714_req_4471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3500_elements(119), ack => phi_stmt_1714_req_0); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(117) & convTransposeA_CP_3500_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1383/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(113) & convTransposeA_CP_3500_elements(116) & convTransposeA_CP_3500_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1383/merge_stmt_1700_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_1383/merge_stmt_1700_PhiAck/$entry
      -- 
    convTransposeA_CP_3500_elements(121) <= OrReduce(convTransposeA_CP_3500_elements(110) & convTransposeA_CP_3500_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1383/merge_stmt_1700_PhiAck/phi_stmt_1701_ack
      -- 
    phi_stmt_1701_ack_4476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1701_ack_0, ack => convTransposeA_CP_3500_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1383/merge_stmt_1700_PhiAck/phi_stmt_1708_ack
      -- 
    phi_stmt_1708_ack_4477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1708_ack_0, ack => convTransposeA_CP_3500_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1383/merge_stmt_1700_PhiAck/phi_stmt_1714_ack
      -- 
    phi_stmt_1714_ack_4478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1714_ack_0, ack => convTransposeA_CP_3500_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1383/merge_stmt_1700_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3500_elements(122) & convTransposeA_CP_3500_elements(123) & convTransposeA_CP_3500_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3500_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1620_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1620_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1597_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1597_scaled : std_logic_vector(13 downto 0);
    signal add41_1451 : std_logic_vector(15 downto 0);
    signal add54_1462 : std_logic_vector(15 downto 0);
    signal add73_1573 : std_logic_vector(63 downto 0);
    signal add75_1583 : std_logic_vector(63 downto 0);
    signal add86_1637 : std_logic_vector(31 downto 0);
    signal add93_1655 : std_logic_vector(15 downto 0);
    signal add_1435 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1531 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1598_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1598_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1598_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1598_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1598_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1598_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1621_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1621_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1621_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1621_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1621_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1621_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1600 : std_logic_vector(31 downto 0);
    signal arrayidx82_1623 : std_logic_vector(31 downto 0);
    signal call11_1404 : std_logic_vector(15 downto 0);
    signal call13_1407 : std_logic_vector(15 downto 0);
    signal call14_1410 : std_logic_vector(15 downto 0);
    signal call15_1413 : std_logic_vector(15 downto 0);
    signal call16_1426 : std_logic_vector(15 downto 0);
    signal call18_1438 : std_logic_vector(15 downto 0);
    signal call1_1389 : std_logic_vector(15 downto 0);
    signal call20_1441 : std_logic_vector(15 downto 0);
    signal call22_1444 : std_logic_vector(15 downto 0);
    signal call3_1392 : std_logic_vector(15 downto 0);
    signal call5_1395 : std_logic_vector(15 downto 0);
    signal call7_1398 : std_logic_vector(15 downto 0);
    signal call9_1401 : std_logic_vector(15 downto 0);
    signal call_1386 : std_logic_vector(15 downto 0);
    signal cmp101_1668 : std_logic_vector(0 downto 0);
    signal cmp112_1693 : std_logic_vector(0 downto 0);
    signal cmp_1642 : std_logic_vector(0 downto 0);
    signal conv107_1688 : std_logic_vector(31 downto 0);
    signal conv110_1483 : std_logic_vector(31 downto 0);
    signal conv17_1430 : std_logic_vector(31 downto 0);
    signal conv61_1555 : std_logic_vector(63 downto 0);
    signal conv64_1471 : std_logic_vector(63 downto 0);
    signal conv66_1559 : std_logic_vector(63 downto 0);
    signal conv69_1475 : std_logic_vector(63 downto 0);
    signal conv71_1563 : std_logic_vector(63 downto 0);
    signal conv85_1631 : std_logic_vector(31 downto 0);
    signal conv89_1479 : std_logic_vector(31 downto 0);
    signal conv_1417 : std_logic_vector(31 downto 0);
    signal idxprom81_1616 : std_logic_vector(63 downto 0);
    signal idxprom_1593 : std_logic_vector(63 downto 0);
    signal inc105_1672 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1677 : std_logic_vector(15 downto 0);
    signal inc_1663 : std_logic_vector(15 downto 0);
    signal indvar_1492 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1726 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1714 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1513 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1708 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1506 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1684 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1701 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1499 : std_logic_vector(15 downto 0);
    signal mul50_1546 : std_logic_vector(15 downto 0);
    signal mul72_1568 : std_logic_vector(63 downto 0);
    signal mul74_1578 : std_logic_vector(63 downto 0);
    signal mul_1536 : std_logic_vector(15 downto 0);
    signal ptr_deref_1603_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1603_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1603_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1603_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1603_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1625_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1625_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1625_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1625_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1625_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1625_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1423 : std_logic_vector(31 downto 0);
    signal shr111126_1489 : std_logic_vector(31 downto 0);
    signal shr80_1610 : std_logic_vector(63 downto 0);
    signal shr_1589 : std_logic_vector(31 downto 0);
    signal sub44_1541 : std_logic_vector(15 downto 0);
    signal sub57_1467 : std_logic_vector(15 downto 0);
    signal sub58_1551 : std_logic_vector(15 downto 0);
    signal sub_1456 : std_logic_vector(15 downto 0);
    signal tmp1_1526 : std_logic_vector(31 downto 0);
    signal tmp78_1604 : std_logic_vector(63 downto 0);
    signal type_cast_1421_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1449_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1460_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1487_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1496_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1498_wire : std_logic_vector(31 downto 0);
    signal type_cast_1503_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1505_wire : std_logic_vector(15 downto 0);
    signal type_cast_1510_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1512_wire : std_logic_vector(15 downto 0);
    signal type_cast_1517_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1519_wire : std_logic_vector(15 downto 0);
    signal type_cast_1524_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1587_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1608_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1614_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1635_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1653_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1661_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1681_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1704_wire : std_logic_vector(15 downto 0);
    signal type_cast_1707_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1711_wire : std_logic_vector(15 downto 0);
    signal type_cast_1713_wire : std_logic_vector(15 downto 0);
    signal type_cast_1717_wire : std_logic_vector(15 downto 0);
    signal type_cast_1719_wire : std_logic_vector(15 downto 0);
    signal type_cast_1724_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1732_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1598_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1598_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1598_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1598_resized_base_address <= "00000000000000";
    array_obj_ref_1621_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1621_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1621_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1621_resized_base_address <= "00000000000000";
    ptr_deref_1603_word_offset_0 <= "00000000000000";
    ptr_deref_1625_word_offset_0 <= "00000000000000";
    type_cast_1421_wire_constant <= "00000000000000000000000000010000";
    type_cast_1449_wire_constant <= "1111111111111111";
    type_cast_1460_wire_constant <= "1111111111111111";
    type_cast_1487_wire_constant <= "00000000000000000000000000000010";
    type_cast_1496_wire_constant <= "00000000000000000000000000000000";
    type_cast_1503_wire_constant <= "0000000000000000";
    type_cast_1510_wire_constant <= "0000000000000000";
    type_cast_1517_wire_constant <= "0000000000000000";
    type_cast_1524_wire_constant <= "00000000000000000000000000000100";
    type_cast_1587_wire_constant <= "00000000000000000000000000000010";
    type_cast_1608_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1614_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1635_wire_constant <= "00000000000000000000000000000100";
    type_cast_1653_wire_constant <= "0000000000000100";
    type_cast_1661_wire_constant <= "0000000000000001";
    type_cast_1681_wire_constant <= "0000000000000000";
    type_cast_1707_wire_constant <= "0000000000000000";
    type_cast_1724_wire_constant <= "00000000000000000000000000000001";
    type_cast_1732_wire_constant <= "0000000000000001";
    phi_stmt_1492: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1496_wire_constant & type_cast_1498_wire;
      req <= phi_stmt_1492_req_0 & phi_stmt_1492_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1492",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1492_ack_0,
          idata => idata,
          odata => indvar_1492,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1492
    phi_stmt_1499: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1503_wire_constant & type_cast_1505_wire;
      req <= phi_stmt_1499_req_0 & phi_stmt_1499_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1499",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1499_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1499,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1499
    phi_stmt_1506: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1510_wire_constant & type_cast_1512_wire;
      req <= phi_stmt_1506_req_0 & phi_stmt_1506_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1506",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1506_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1506,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1506
    phi_stmt_1513: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1517_wire_constant & type_cast_1519_wire;
      req <= phi_stmt_1513_req_0 & phi_stmt_1513_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1513",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1513_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1513,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1513
    phi_stmt_1701: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1704_wire & type_cast_1707_wire_constant;
      req <= phi_stmt_1701_req_0 & phi_stmt_1701_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1701",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1701_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1701,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1701
    phi_stmt_1708: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1711_wire & type_cast_1713_wire;
      req <= phi_stmt_1708_req_0 & phi_stmt_1708_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1708",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1708_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1708,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1708
    phi_stmt_1714: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1717_wire & type_cast_1719_wire;
      req <= phi_stmt_1714_req_0 & phi_stmt_1714_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1714",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1714_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1714,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1714
    -- flow-through select operator MUX_1683_inst
    input_dim1x_x2_1684 <= type_cast_1681_wire_constant when (cmp101_1668(0) /=  '0') else inc_1663;
    addr_of_1599_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1599_final_reg_req_0;
      addr_of_1599_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1599_final_reg_req_1;
      addr_of_1599_final_reg_ack_1<= rack(0);
      addr_of_1599_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1599_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1598_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1622_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1622_final_reg_req_0;
      addr_of_1622_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1622_final_reg_req_1;
      addr_of_1622_final_reg_ack_1<= rack(0);
      addr_of_1622_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1622_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1621_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1623,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1416_inst_req_0;
      type_cast_1416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1416_inst_req_1;
      type_cast_1416_inst_ack_1<= rack(0);
      type_cast_1416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1429_inst_req_0;
      type_cast_1429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1429_inst_req_1;
      type_cast_1429_inst_ack_1<= rack(0);
      type_cast_1429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1430,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1470_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1470_inst_req_0;
      type_cast_1470_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1470_inst_req_1;
      type_cast_1470_inst_ack_1<= rack(0);
      type_cast_1470_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1470_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1471,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1474_inst_req_0;
      type_cast_1474_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1474_inst_req_1;
      type_cast_1474_inst_ack_1<= rack(0);
      type_cast_1474_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1474_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1478_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1478_inst_req_0;
      type_cast_1478_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1478_inst_req_1;
      type_cast_1478_inst_ack_1<= rack(0);
      type_cast_1478_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1478_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1482_inst_req_0;
      type_cast_1482_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1482_inst_req_1;
      type_cast_1482_inst_ack_1<= rack(0);
      type_cast_1482_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1482_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1498_inst_req_0;
      type_cast_1498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1498_inst_req_1;
      type_cast_1498_inst_ack_1<= rack(0);
      type_cast_1498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1498_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1505_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1505_inst_req_0;
      type_cast_1505_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1505_inst_req_1;
      type_cast_1505_inst_ack_1<= rack(0);
      type_cast_1505_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1505_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1701,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1505_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1512_inst_req_0;
      type_cast_1512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1512_inst_req_1;
      type_cast_1512_inst_ack_1<= rack(0);
      type_cast_1512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1512_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1519_inst_req_0;
      type_cast_1519_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1519_inst_req_1;
      type_cast_1519_inst_ack_1<= rack(0);
      type_cast_1519_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1519_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1519_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1554_inst_req_0;
      type_cast_1554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1554_inst_req_1;
      type_cast_1554_inst_ack_1<= rack(0);
      type_cast_1554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1555,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1558_inst_req_0;
      type_cast_1558_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1558_inst_req_1;
      type_cast_1558_inst_ack_1<= rack(0);
      type_cast_1558_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1558_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1559,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1562_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1562_inst_req_0;
      type_cast_1562_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1562_inst_req_1;
      type_cast_1562_inst_ack_1<= rack(0);
      type_cast_1562_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1562_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1563,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1592_inst_req_0;
      type_cast_1592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1592_inst_req_1;
      type_cast_1592_inst_ack_1<= rack(0);
      type_cast_1592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1630_inst_req_0;
      type_cast_1630_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1630_inst_req_1;
      type_cast_1630_inst_ack_1<= rack(0);
      type_cast_1630_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1630_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1671_inst_req_0;
      type_cast_1671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1671_inst_req_1;
      type_cast_1671_inst_ack_1<= rack(0);
      type_cast_1671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1668,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1687_inst_req_0;
      type_cast_1687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1687_inst_req_1;
      type_cast_1687_inst_ack_1<= rack(0);
      type_cast_1687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1677,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1704_inst_req_0;
      type_cast_1704_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1704_inst_req_1;
      type_cast_1704_inst_ack_1<= rack(0);
      type_cast_1704_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1704_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1704_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1711_inst_req_0;
      type_cast_1711_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1711_inst_req_1;
      type_cast_1711_inst_ack_1<= rack(0);
      type_cast_1711_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1711_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1713_inst_req_0;
      type_cast_1713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1713_inst_req_1;
      type_cast_1713_inst_ack_1<= rack(0);
      type_cast_1713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1713_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1717_inst_req_0;
      type_cast_1717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1717_inst_req_1;
      type_cast_1717_inst_ack_1<= rack(0);
      type_cast_1717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1717_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1513,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1717_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1719_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1719_inst_req_0;
      type_cast_1719_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1719_inst_req_1;
      type_cast_1719_inst_ack_1<= rack(0);
      type_cast_1719_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1719_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1677,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1719_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1598_index_1_rename
    process(R_idxprom_1597_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1597_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1597_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1598_index_1_resize
    process(idxprom_1593) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1593;
      ov := iv(13 downto 0);
      R_idxprom_1597_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1598_root_address_inst
    process(array_obj_ref_1598_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1598_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1598_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1621_index_1_rename
    process(R_idxprom81_1620_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1620_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1620_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1621_index_1_resize
    process(idxprom81_1616) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1616;
      ov := iv(13 downto 0);
      R_idxprom81_1620_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1621_root_address_inst
    process(array_obj_ref_1621_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1621_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1621_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1603_addr_0
    process(ptr_deref_1603_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1603_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1603_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1603_base_resize
    process(arrayidx77_1600) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1600;
      ov := iv(13 downto 0);
      ptr_deref_1603_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1603_gather_scatter
    process(ptr_deref_1603_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1603_data_0;
      ov(63 downto 0) := iv;
      tmp78_1604 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1603_root_address_inst
    process(ptr_deref_1603_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1603_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1603_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1625_addr_0
    process(ptr_deref_1625_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1625_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1625_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1625_base_resize
    process(arrayidx82_1623) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1623;
      ov := iv(13 downto 0);
      ptr_deref_1625_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1625_gather_scatter
    process(tmp78_1604) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1604;
      ov(63 downto 0) := iv;
      ptr_deref_1625_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1625_root_address_inst
    process(ptr_deref_1625_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1625_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1625_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1643_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1642;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1643_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1643_branch_req_0,
          ack0 => if_stmt_1643_branch_ack_0,
          ack1 => if_stmt_1643_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1694_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1693;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1694_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1694_branch_req_0,
          ack0 => if_stmt_1694_branch_ack_0,
          ack1 => if_stmt_1694_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1450_inst
    process(call7_1398) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1398, type_cast_1449_wire_constant, tmp_var);
      add41_1451 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1461_inst
    process(call9_1401) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1401, type_cast_1460_wire_constant, tmp_var);
      add54_1462 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1540_inst
    process(sub_1456, mul_1536) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1456, mul_1536, tmp_var);
      sub44_1541 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1550_inst
    process(sub57_1467, mul50_1546) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1467, mul50_1546, tmp_var);
      sub58_1551 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1654_inst
    process(input_dim2x_x1_1499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1499, type_cast_1653_wire_constant, tmp_var);
      add93_1655 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1662_inst
    process(input_dim1x_x1_1506) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1506, type_cast_1661_wire_constant, tmp_var);
      inc_1663 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1676_inst
    process(inc105_1672, input_dim0x_x2_1513) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1672, input_dim0x_x2_1513, tmp_var);
      inc105x_xinput_dim0x_x2_1677 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1530_inst
    process(add_1435, tmp1_1526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1435, tmp1_1526, tmp_var);
      add_src_0x_x0_1531 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1636_inst
    process(conv85_1631) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1631, type_cast_1635_wire_constant, tmp_var);
      add86_1637 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1725_inst
    process(indvar_1492) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1492, type_cast_1724_wire_constant, tmp_var);
      indvarx_xnext_1726 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1572_inst
    process(mul72_1568, conv66_1559) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1568, conv66_1559, tmp_var);
      add73_1573 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1582_inst
    process(mul74_1578, conv61_1555) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1578, conv61_1555, tmp_var);
      add75_1583 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1615_inst
    process(shr80_1610) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1610, type_cast_1614_wire_constant, tmp_var);
      idxprom81_1616 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1667_inst
    process(inc_1663, call1_1389) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1663, call1_1389, tmp_var);
      cmp101_1668 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1692_inst
    process(conv107_1688, shr111126_1489) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1688, shr111126_1489, tmp_var);
      cmp112_1693 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1488_inst
    process(conv110_1483) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1483, type_cast_1487_wire_constant, tmp_var);
      shr111126_1489 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1588_inst
    process(add_src_0x_x0_1531) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1531, type_cast_1587_wire_constant, tmp_var);
      shr_1589 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1609_inst
    process(add75_1583) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1583, type_cast_1608_wire_constant, tmp_var);
      shr80_1610 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1535_inst
    process(input_dim0x_x2_1513, call13_1407) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1513, call13_1407, tmp_var);
      mul_1536 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1545_inst
    process(input_dim1x_x1_1506, call13_1407) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1506, call13_1407, tmp_var);
      mul50_1546 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1525_inst
    process(indvar_1492) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1492, type_cast_1524_wire_constant, tmp_var);
      tmp1_1526 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1567_inst
    process(conv71_1563, conv69_1475) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1563, conv69_1475, tmp_var);
      mul72_1568 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1577_inst
    process(add73_1573, conv64_1471) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1573, conv64_1471, tmp_var);
      mul74_1578 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1434_inst
    process(shl_1423, conv17_1430) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1423, conv17_1430, tmp_var);
      add_1435 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1422_inst
    process(conv_1417) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1417, type_cast_1421_wire_constant, tmp_var);
      shl_1423 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1455_inst
    process(add41_1451, call14_1410) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1451, call14_1410, tmp_var);
      sub_1456 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1466_inst
    process(add54_1462, call14_1410) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1462, call14_1410, tmp_var);
      sub57_1467 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1641_inst
    process(add86_1637, conv89_1479) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1637, conv89_1479, tmp_var);
      cmp_1642 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1598_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1597_scaled;
      array_obj_ref_1598_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1598_index_offset_req_0;
      array_obj_ref_1598_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1598_index_offset_req_1;
      array_obj_ref_1598_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1621_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1620_scaled;
      array_obj_ref_1621_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1621_index_offset_req_0;
      array_obj_ref_1621_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1621_index_offset_req_1;
      array_obj_ref_1621_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1603_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1603_load_0_req_0;
      ptr_deref_1603_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1603_load_0_req_1;
      ptr_deref_1603_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1603_word_address_0;
      ptr_deref_1603_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1625_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1625_store_0_req_0;
      ptr_deref_1625_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1625_store_0_req_1;
      ptr_deref_1625_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1625_word_address_0;
      data_in <= ptr_deref_1625_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1385_inst RPIPE_Block0_start_1388_inst RPIPE_Block0_start_1391_inst RPIPE_Block0_start_1394_inst RPIPE_Block0_start_1397_inst RPIPE_Block0_start_1400_inst RPIPE_Block0_start_1403_inst RPIPE_Block0_start_1406_inst RPIPE_Block0_start_1409_inst RPIPE_Block0_start_1412_inst RPIPE_Block0_start_1425_inst RPIPE_Block0_start_1437_inst RPIPE_Block0_start_1440_inst RPIPE_Block0_start_1443_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1385_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1388_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1391_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1394_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1397_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1400_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1403_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1406_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1409_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1412_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1425_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1437_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1440_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1443_inst_req_0;
      RPIPE_Block0_start_1385_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1388_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1391_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1394_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1397_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1400_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1403_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1406_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1409_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1412_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1425_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1437_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1440_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1443_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1385_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1388_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1391_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1394_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1397_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1400_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1403_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1406_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1409_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1412_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1425_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1437_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1440_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1443_inst_req_1;
      RPIPE_Block0_start_1385_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1388_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1391_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1394_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1397_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1400_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1403_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1406_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1409_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1412_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1425_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1437_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1440_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1443_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_1386 <= data_out(223 downto 208);
      call1_1389 <= data_out(207 downto 192);
      call3_1392 <= data_out(191 downto 176);
      call5_1395 <= data_out(175 downto 160);
      call7_1398 <= data_out(159 downto 144);
      call9_1401 <= data_out(143 downto 128);
      call11_1404 <= data_out(127 downto 112);
      call13_1407 <= data_out(111 downto 96);
      call14_1410 <= data_out(95 downto 80);
      call15_1413 <= data_out(79 downto 64);
      call16_1426 <= data_out(63 downto 48);
      call18_1438 <= data_out(47 downto 32);
      call20_1441 <= data_out(31 downto 16);
      call22_1444 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1730_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1730_inst_req_0;
      WPIPE_Block0_done_1730_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1730_inst_req_1;
      WPIPE_Block0_done_1730_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1732_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4495_start: Boolean;
  signal convTransposeB_CP_4495_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2032_inst_req_0 : boolean;
  signal ptr_deref_1986_store_0_ack_1 : boolean;
  signal ptr_deref_1986_store_0_req_1 : boolean;
  signal addr_of_1960_final_reg_ack_1 : boolean;
  signal type_cast_2032_inst_ack_0 : boolean;
  signal addr_of_1960_final_reg_req_1 : boolean;
  signal type_cast_1991_inst_req_0 : boolean;
  signal type_cast_1991_inst_ack_0 : boolean;
  signal array_obj_ref_1959_index_offset_req_0 : boolean;
  signal if_stmt_2004_branch_req_0 : boolean;
  signal if_stmt_2004_branch_ack_1 : boolean;
  signal addr_of_1983_final_reg_req_0 : boolean;
  signal type_cast_1991_inst_ack_1 : boolean;
  signal addr_of_1983_final_reg_ack_0 : boolean;
  signal RPIPE_Block1_start_1741_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1741_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1741_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1741_inst_ack_1 : boolean;
  signal addr_of_1960_final_reg_ack_0 : boolean;
  signal addr_of_1983_final_reg_req_1 : boolean;
  signal addr_of_1983_final_reg_ack_1 : boolean;
  signal WPIPE_Block1_done_2091_inst_req_0 : boolean;
  signal ptr_deref_1964_load_0_req_0 : boolean;
  signal WPIPE_Block1_done_2091_inst_ack_0 : boolean;
  signal ptr_deref_1964_load_0_ack_0 : boolean;
  signal type_cast_1880_inst_req_0 : boolean;
  signal array_obj_ref_1959_index_offset_ack_0 : boolean;
  signal type_cast_1880_inst_req_1 : boolean;
  signal type_cast_1880_inst_ack_0 : boolean;
  signal if_stmt_2004_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2091_inst_req_1 : boolean;
  signal type_cast_1991_inst_req_1 : boolean;
  signal ptr_deref_1964_load_0_req_1 : boolean;
  signal WPIPE_Block1_done_2091_inst_ack_1 : boolean;
  signal ptr_deref_1964_load_0_ack_1 : boolean;
  signal type_cast_1880_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1744_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1744_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1744_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1744_inst_ack_1 : boolean;
  signal if_stmt_2055_branch_ack_0 : boolean;
  signal RPIPE_Block1_start_1747_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1747_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1747_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1747_inst_ack_1 : boolean;
  signal if_stmt_2055_branch_ack_1 : boolean;
  signal array_obj_ref_1982_index_offset_ack_1 : boolean;
  signal RPIPE_Block1_start_1750_inst_req_0 : boolean;
  signal ptr_deref_1986_store_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1750_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1750_inst_req_1 : boolean;
  signal ptr_deref_1986_store_0_req_0 : boolean;
  signal RPIPE_Block1_start_1750_inst_ack_1 : boolean;
  signal if_stmt_2055_branch_req_0 : boolean;
  signal array_obj_ref_1982_index_offset_req_1 : boolean;
  signal RPIPE_Block1_start_1753_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1753_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1753_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1753_inst_ack_1 : boolean;
  signal type_cast_2048_inst_ack_1 : boolean;
  signal array_obj_ref_1982_index_offset_ack_0 : boolean;
  signal array_obj_ref_1982_index_offset_req_0 : boolean;
  signal RPIPE_Block1_start_1756_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1756_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1756_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1756_inst_ack_1 : boolean;
  signal addr_of_1960_final_reg_req_0 : boolean;
  signal RPIPE_Block1_start_1759_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1759_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1759_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1759_inst_ack_1 : boolean;
  signal array_obj_ref_1959_index_offset_ack_1 : boolean;
  signal array_obj_ref_1959_index_offset_req_1 : boolean;
  signal type_cast_2048_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1762_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1762_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1762_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1762_inst_ack_1 : boolean;
  signal type_cast_2048_inst_ack_0 : boolean;
  signal type_cast_2048_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1765_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1765_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1765_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1765_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1768_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1768_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1768_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1768_inst_ack_1 : boolean;
  signal type_cast_2032_inst_ack_1 : boolean;
  signal type_cast_2032_inst_req_1 : boolean;
  signal type_cast_1772_inst_req_0 : boolean;
  signal type_cast_1772_inst_ack_0 : boolean;
  signal type_cast_1772_inst_req_1 : boolean;
  signal type_cast_1772_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1781_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1781_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1781_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1781_inst_ack_1 : boolean;
  signal type_cast_1785_inst_req_0 : boolean;
  signal type_cast_1785_inst_ack_0 : boolean;
  signal type_cast_1785_inst_req_1 : boolean;
  signal type_cast_1785_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1793_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1793_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1793_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1793_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1796_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1796_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1796_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1796_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1799_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1799_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1799_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1799_inst_ack_1 : boolean;
  signal type_cast_1832_inst_req_0 : boolean;
  signal type_cast_1832_inst_ack_0 : boolean;
  signal type_cast_1832_inst_req_1 : boolean;
  signal type_cast_1832_inst_ack_1 : boolean;
  signal type_cast_1836_inst_req_0 : boolean;
  signal type_cast_1836_inst_ack_0 : boolean;
  signal type_cast_1836_inst_req_1 : boolean;
  signal type_cast_1836_inst_ack_1 : boolean;
  signal type_cast_1840_inst_req_0 : boolean;
  signal type_cast_1840_inst_ack_0 : boolean;
  signal type_cast_1840_inst_req_1 : boolean;
  signal type_cast_1840_inst_ack_1 : boolean;
  signal type_cast_1844_inst_req_0 : boolean;
  signal type_cast_1844_inst_ack_0 : boolean;
  signal type_cast_1844_inst_req_1 : boolean;
  signal type_cast_1844_inst_ack_1 : boolean;
  signal type_cast_1915_inst_req_0 : boolean;
  signal type_cast_1915_inst_ack_0 : boolean;
  signal type_cast_1915_inst_req_1 : boolean;
  signal type_cast_1915_inst_ack_1 : boolean;
  signal type_cast_1919_inst_req_0 : boolean;
  signal type_cast_1919_inst_ack_0 : boolean;
  signal type_cast_1919_inst_req_1 : boolean;
  signal type_cast_1919_inst_ack_1 : boolean;
  signal type_cast_1923_inst_req_0 : boolean;
  signal type_cast_1923_inst_ack_0 : boolean;
  signal type_cast_1923_inst_req_1 : boolean;
  signal type_cast_1923_inst_ack_1 : boolean;
  signal type_cast_1953_inst_req_0 : boolean;
  signal type_cast_1953_inst_ack_0 : boolean;
  signal type_cast_1953_inst_req_1 : boolean;
  signal type_cast_1953_inst_ack_1 : boolean;
  signal phi_stmt_1875_req_1 : boolean;
  signal phi_stmt_1868_req_0 : boolean;
  signal phi_stmt_1861_req_0 : boolean;
  signal phi_stmt_1854_req_1 : boolean;
  signal type_cast_1878_inst_req_0 : boolean;
  signal type_cast_1878_inst_ack_0 : boolean;
  signal type_cast_1878_inst_req_1 : boolean;
  signal type_cast_1878_inst_ack_1 : boolean;
  signal phi_stmt_1875_req_0 : boolean;
  signal type_cast_1874_inst_req_0 : boolean;
  signal type_cast_1874_inst_ack_0 : boolean;
  signal type_cast_1874_inst_req_1 : boolean;
  signal type_cast_1874_inst_ack_1 : boolean;
  signal phi_stmt_1868_req_1 : boolean;
  signal type_cast_1867_inst_req_0 : boolean;
  signal type_cast_1867_inst_ack_0 : boolean;
  signal type_cast_1867_inst_req_1 : boolean;
  signal type_cast_1867_inst_ack_1 : boolean;
  signal phi_stmt_1861_req_1 : boolean;
  signal type_cast_1857_inst_req_0 : boolean;
  signal type_cast_1857_inst_ack_0 : boolean;
  signal type_cast_1857_inst_req_1 : boolean;
  signal type_cast_1857_inst_ack_1 : boolean;
  signal phi_stmt_1854_req_0 : boolean;
  signal phi_stmt_1854_ack_0 : boolean;
  signal phi_stmt_1861_ack_0 : boolean;
  signal phi_stmt_1868_ack_0 : boolean;
  signal phi_stmt_1875_ack_0 : boolean;
  signal type_cast_2080_inst_req_0 : boolean;
  signal type_cast_2080_inst_ack_0 : boolean;
  signal type_cast_2080_inst_req_1 : boolean;
  signal type_cast_2080_inst_ack_1 : boolean;
  signal phi_stmt_2075_req_1 : boolean;
  signal type_cast_2074_inst_req_0 : boolean;
  signal type_cast_2074_inst_ack_0 : boolean;
  signal type_cast_2074_inst_req_1 : boolean;
  signal type_cast_2074_inst_ack_1 : boolean;
  signal phi_stmt_2069_req_1 : boolean;
  signal phi_stmt_2062_req_1 : boolean;
  signal type_cast_2078_inst_req_0 : boolean;
  signal type_cast_2078_inst_ack_0 : boolean;
  signal type_cast_2078_inst_req_1 : boolean;
  signal type_cast_2078_inst_ack_1 : boolean;
  signal phi_stmt_2075_req_0 : boolean;
  signal type_cast_2072_inst_req_0 : boolean;
  signal type_cast_2072_inst_ack_0 : boolean;
  signal type_cast_2072_inst_req_1 : boolean;
  signal type_cast_2072_inst_ack_1 : boolean;
  signal phi_stmt_2069_req_0 : boolean;
  signal type_cast_2065_inst_req_0 : boolean;
  signal type_cast_2065_inst_ack_0 : boolean;
  signal type_cast_2065_inst_req_1 : boolean;
  signal type_cast_2065_inst_ack_1 : boolean;
  signal phi_stmt_2062_req_0 : boolean;
  signal phi_stmt_2062_ack_0 : boolean;
  signal phi_stmt_2069_ack_0 : boolean;
  signal phi_stmt_2075_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4495_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4495_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4495_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4495_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4495: Block -- control-path 
    signal convTransposeB_CP_4495_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4495_elements(0) <= convTransposeB_CP_4495_start;
    convTransposeB_CP_4495_symbol <= convTransposeB_CP_4495_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/branch_block_stmt_1739__entry__
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800__entry__
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Update/cr
      -- 
    rr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(0), ack => RPIPE_Block1_start_1741_inst_req_0); -- 
    cr_4688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(0), ack => type_cast_1772_inst_req_1); -- 
    cr_4716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(0), ack => type_cast_1785_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1739/assign_stmt_2087__exit__
      -- CP-element group 1: 	 branch_block_stmt_1739/assign_stmt_2087__entry__
      -- CP-element group 1: 	 branch_block_stmt_1739/merge_stmt_2061__exit__
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1739/assign_stmt_2087/$exit
      -- CP-element group 1: 	 branch_block_stmt_1739/assign_stmt_2087/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/cr
      -- 
    rr_5244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1878_inst_req_0); -- 
    cr_5249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1878_inst_req_1); -- 
    rr_5267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1874_inst_req_0); -- 
    cr_5272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1874_inst_req_1); -- 
    rr_5290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1867_inst_req_0); -- 
    cr_5295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1867_inst_req_1); -- 
    rr_5313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1857_inst_req_0); -- 
    cr_5318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(1), ack => type_cast_1857_inst_req_1); -- 
    convTransposeB_CP_4495_elements(1) <= convTransposeB_CP_4495_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Update/cr
      -- 
    ra_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1741_inst_ack_0, ack => convTransposeB_CP_4495_elements(2)); -- 
    cr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(2), ack => RPIPE_Block1_start_1741_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1741_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Sample/rr
      -- 
    ca_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1741_inst_ack_1, ack => convTransposeB_CP_4495_elements(3)); -- 
    rr_4557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(3), ack => RPIPE_Block1_start_1744_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Update/cr
      -- 
    ra_4558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1744_inst_ack_0, ack => convTransposeB_CP_4495_elements(4)); -- 
    cr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(4), ack => RPIPE_Block1_start_1744_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1744_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Sample/rr
      -- 
    ca_4563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1744_inst_ack_1, ack => convTransposeB_CP_4495_elements(5)); -- 
    rr_4571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(5), ack => RPIPE_Block1_start_1747_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Update/cr
      -- 
    ra_4572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1747_inst_ack_0, ack => convTransposeB_CP_4495_elements(6)); -- 
    cr_4576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(6), ack => RPIPE_Block1_start_1747_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1747_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Sample/rr
      -- 
    ca_4577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1747_inst_ack_1, ack => convTransposeB_CP_4495_elements(7)); -- 
    rr_4585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(7), ack => RPIPE_Block1_start_1750_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Update/cr
      -- 
    ra_4586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1750_inst_ack_0, ack => convTransposeB_CP_4495_elements(8)); -- 
    cr_4590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(8), ack => RPIPE_Block1_start_1750_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1750_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Sample/rr
      -- 
    ca_4591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1750_inst_ack_1, ack => convTransposeB_CP_4495_elements(9)); -- 
    rr_4599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(9), ack => RPIPE_Block1_start_1753_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Update/cr
      -- 
    ra_4600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1753_inst_ack_0, ack => convTransposeB_CP_4495_elements(10)); -- 
    cr_4604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(10), ack => RPIPE_Block1_start_1753_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1753_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Sample/rr
      -- 
    ca_4605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1753_inst_ack_1, ack => convTransposeB_CP_4495_elements(11)); -- 
    rr_4613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(11), ack => RPIPE_Block1_start_1756_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Update/cr
      -- 
    ra_4614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1756_inst_ack_0, ack => convTransposeB_CP_4495_elements(12)); -- 
    cr_4618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(12), ack => RPIPE_Block1_start_1756_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1756_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Sample/rr
      -- 
    ca_4619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1756_inst_ack_1, ack => convTransposeB_CP_4495_elements(13)); -- 
    rr_4627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(13), ack => RPIPE_Block1_start_1759_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Update/cr
      -- 
    ra_4628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1759_inst_ack_0, ack => convTransposeB_CP_4495_elements(14)); -- 
    cr_4632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(14), ack => RPIPE_Block1_start_1759_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1759_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Sample/rr
      -- 
    ca_4633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1759_inst_ack_1, ack => convTransposeB_CP_4495_elements(15)); -- 
    rr_4641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(15), ack => RPIPE_Block1_start_1762_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Update/cr
      -- 
    ra_4642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1762_inst_ack_0, ack => convTransposeB_CP_4495_elements(16)); -- 
    cr_4646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(16), ack => RPIPE_Block1_start_1762_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1762_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Sample/rr
      -- 
    ca_4647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1762_inst_ack_1, ack => convTransposeB_CP_4495_elements(17)); -- 
    rr_4655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(17), ack => RPIPE_Block1_start_1765_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Update/cr
      -- 
    ra_4656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1765_inst_ack_0, ack => convTransposeB_CP_4495_elements(18)); -- 
    cr_4660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(18), ack => RPIPE_Block1_start_1765_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1765_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Sample/rr
      -- 
    ca_4661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1765_inst_ack_1, ack => convTransposeB_CP_4495_elements(19)); -- 
    rr_4669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(19), ack => RPIPE_Block1_start_1768_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Update/cr
      -- 
    ra_4670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1768_inst_ack_0, ack => convTransposeB_CP_4495_elements(20)); -- 
    cr_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(20), ack => RPIPE_Block1_start_1768_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1768_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Sample/rr
      -- 
    ca_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1768_inst_ack_1, ack => convTransposeB_CP_4495_elements(21)); -- 
    rr_4683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(21), ack => type_cast_1772_inst_req_0); -- 
    rr_4697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(21), ack => RPIPE_Block1_start_1781_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Sample/ra
      -- 
    ra_4684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_0, ack => convTransposeB_CP_4495_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1772_Update/ca
      -- 
    ca_4689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_1, ack => convTransposeB_CP_4495_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Update/cr
      -- 
    ra_4698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1781_inst_ack_0, ack => convTransposeB_CP_4495_elements(24)); -- 
    cr_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(24), ack => RPIPE_Block1_start_1781_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1781_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Sample/rr
      -- 
    ca_4703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1781_inst_ack_1, ack => convTransposeB_CP_4495_elements(25)); -- 
    rr_4711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(25), ack => type_cast_1785_inst_req_0); -- 
    rr_4725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(25), ack => RPIPE_Block1_start_1793_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Sample/ra
      -- 
    ra_4712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_0, ack => convTransposeB_CP_4495_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/type_cast_1785_Update/ca
      -- 
    ca_4717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_1, ack => convTransposeB_CP_4495_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Update/cr
      -- 
    ra_4726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1793_inst_ack_0, ack => convTransposeB_CP_4495_elements(28)); -- 
    cr_4730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(28), ack => RPIPE_Block1_start_1793_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1793_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Sample/rr
      -- 
    ca_4731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1793_inst_ack_1, ack => convTransposeB_CP_4495_elements(29)); -- 
    rr_4739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(29), ack => RPIPE_Block1_start_1796_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Update/cr
      -- 
    ra_4740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1796_inst_ack_0, ack => convTransposeB_CP_4495_elements(30)); -- 
    cr_4744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(30), ack => RPIPE_Block1_start_1796_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1796_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Sample/rr
      -- 
    ca_4745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1796_inst_ack_1, ack => convTransposeB_CP_4495_elements(31)); -- 
    rr_4753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(31), ack => RPIPE_Block1_start_1799_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Update/cr
      -- 
    ra_4754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1799_inst_ack_0, ack => convTransposeB_CP_4495_elements(32)); -- 
    cr_4758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(32), ack => RPIPE_Block1_start_1799_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/RPIPE_Block1_start_1799_Update/ca
      -- 
    ca_4759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1799_inst_ack_1, ack => convTransposeB_CP_4495_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800/$exit
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851__entry__
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1742_to_assign_stmt_1800__exit__
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Update/cr
      -- 
    rr_4770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1832_inst_req_0); -- 
    cr_4775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1832_inst_req_1); -- 
    rr_4784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1836_inst_req_0); -- 
    cr_4789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1836_inst_req_1); -- 
    rr_4798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1840_inst_req_0); -- 
    cr_4803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1840_inst_req_1); -- 
    rr_4812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1844_inst_req_0); -- 
    cr_4817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(34), ack => type_cast_1844_inst_req_1); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(23) & convTransposeB_CP_4495_elements(27) & convTransposeB_CP_4495_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Sample/ra
      -- 
    ra_4771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_0, ack => convTransposeB_CP_4495_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1832_Update/ca
      -- 
    ca_4776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_1, ack => convTransposeB_CP_4495_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Sample/ra
      -- 
    ra_4785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1836_inst_ack_0, ack => convTransposeB_CP_4495_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1836_Update/ca
      -- 
    ca_4790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1836_inst_ack_1, ack => convTransposeB_CP_4495_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Sample/ra
      -- 
    ra_4799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1840_inst_ack_0, ack => convTransposeB_CP_4495_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1840_Update/ca
      -- 
    ca_4804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1840_inst_ack_1, ack => convTransposeB_CP_4495_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Sample/ra
      -- 
    ra_4813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1844_inst_ack_0, ack => convTransposeB_CP_4495_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/type_cast_1844_Update/ca
      -- 
    ca_4818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1844_inst_ack_1, ack => convTransposeB_CP_4495_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851__exit__
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/assign_stmt_1807_to_assign_stmt_1851/$exit
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1868/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1861/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1854/$entry
      -- CP-element group 43: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$entry
      -- 
    rr_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(43), ack => type_cast_1880_inst_req_0); -- 
    cr_5199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(43), ack => type_cast_1880_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(36) & convTransposeB_CP_4495_elements(38) & convTransposeB_CP_4495_elements(40) & convTransposeB_CP_4495_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Sample/ra
      -- 
    ra_4830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1915_inst_ack_0, ack => convTransposeB_CP_4495_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Update/ca
      -- 
    ca_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1915_inst_ack_1, ack => convTransposeB_CP_4495_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Sample/ra
      -- 
    ra_4844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_0, ack => convTransposeB_CP_4495_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Update/ca
      -- 
    ca_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_1, ack => convTransposeB_CP_4495_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Sample/ra
      -- 
    ra_4858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_0, ack => convTransposeB_CP_4495_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Update/ca
      -- 
    ca_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_1, ack => convTransposeB_CP_4495_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Sample/ra
      -- 
    ra_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_0, ack => convTransposeB_CP_4495_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_index_scale_1/scale_rename_req
      -- 
    ca_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_1, ack => convTransposeB_CP_4495_elements(51)); -- 
    req_4902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(51), ack => array_obj_ref_1959_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Sample/ack
      -- 
    ack_4903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1959_index_offset_ack_0, ack => convTransposeB_CP_4495_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_request/req
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_offset_calculated
      -- 
    ack_4908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1959_index_offset_ack_1, ack => convTransposeB_CP_4495_elements(53)); -- 
    req_4917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(53), ack => addr_of_1960_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_request/ack
      -- CP-element group 54: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_sample_completed_
      -- 
    ack_4918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1960_final_reg_ack_0, ack => convTransposeB_CP_4495_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/word_access_start/word_0/rr
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_update_completed_
      -- 
    ack_4923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1960_final_reg_ack_1, ack => convTransposeB_CP_4495_elements(55)); -- 
    rr_4956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(55), ack => ptr_deref_1964_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Sample/word_access_start/word_0/ra
      -- 
    ra_4957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_load_0_ack_0, ack => convTransposeB_CP_4495_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/ptr_deref_1964_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/ptr_deref_1964_Merge/merge_ack
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/ptr_deref_1964_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/ptr_deref_1964_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_update_completed_
      -- 
    ca_4968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_load_0_ack_1, ack => convTransposeB_CP_4495_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_index_scaled_1
      -- 
    req_4998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(58), ack => array_obj_ref_1982_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(45) & convTransposeB_CP_4495_elements(47) & convTransposeB_CP_4495_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_sample_complete
      -- 
    ack_4999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1982_index_offset_ack_0, ack => convTransposeB_CP_4495_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_request/req
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Update/$exit
      -- 
    ack_5004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1982_index_offset_ack_1, ack => convTransposeB_CP_4495_elements(60)); -- 
    req_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(60), ack => addr_of_1983_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_request/ack
      -- CP-element group 61: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_request/$exit
      -- 
    ack_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1983_final_reg_ack_0, ack => convTransposeB_CP_4495_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_word_addrgen/root_register_req
      -- 
    ack_5019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1983_final_reg_ack_1, ack => convTransposeB_CP_4495_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/word_access_start/word_0/rr
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/ptr_deref_1986_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/ptr_deref_1986_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/ptr_deref_1986_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/ptr_deref_1986_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/$entry
      -- 
    rr_5057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(63), ack => ptr_deref_1986_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(57) & convTransposeB_CP_4495_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/word_access_start/word_0/ra
      -- CP-element group 64: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Sample/$exit
      -- 
    ra_5058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1986_store_0_ack_0, ack => convTransposeB_CP_4495_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/word_access_complete/word_0/ca
      -- CP-element group 65: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/$exit
      -- 
    ca_5069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1986_store_0_ack_1, ack => convTransposeB_CP_4495_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Sample/ra
      -- 
    ra_5078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1991_inst_ack_0, ack => convTransposeB_CP_4495_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Update/$exit
      -- 
    ca_5083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1991_inst_ack_1, ack => convTransposeB_CP_4495_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1739/if_stmt_2004_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1739/if_stmt_2004_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1739/if_stmt_2004_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1739/if_stmt_2004_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1739/if_stmt_2004_else_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1739/R_cmp_2005_place
      -- CP-element group 68: 	 branch_block_stmt_1739/if_stmt_2004_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1739/if_stmt_2004__entry__
      -- CP-element group 68: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003__exit__
      -- CP-element group 68: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/$exit
      -- 
    branch_req_5091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(68), ack => if_stmt_2004_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(52) & convTransposeB_CP_4495_elements(59) & convTransposeB_CP_4495_elements(65) & convTransposeB_CP_4495_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1739/merge_stmt_2010_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1739/assign_stmt_2016/$exit
      -- CP-element group 69: 	 branch_block_stmt_1739/assign_stmt_2016/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/if_stmt_2004_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1739/if_stmt_2004_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1739/assign_stmt_2016__exit__
      -- CP-element group 69: 	 branch_block_stmt_1739/assign_stmt_2016__entry__
      -- CP-element group 69: 	 branch_block_stmt_1739/merge_stmt_2010__exit__
      -- CP-element group 69: 	 branch_block_stmt_1739/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1739/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1739/merge_stmt_2010_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/merge_stmt_2010_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1739/merge_stmt_2010_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2004_branch_ack_1, ack => convTransposeB_CP_4495_elements(69)); -- 
    rr_5428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(69), ack => type_cast_2078_inst_req_0); -- 
    cr_5433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(69), ack => type_cast_2078_inst_req_1); -- 
    rr_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(69), ack => type_cast_2072_inst_req_0); -- 
    cr_5456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(69), ack => type_cast_2072_inst_req_1); -- 
    rr_5474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(69), ack => type_cast_2065_inst_req_0); -- 
    cr_5479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(69), ack => type_cast_2065_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1739/merge_stmt_2018_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/$entry
      -- CP-element group 70: 	 branch_block_stmt_1739/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1739/if_stmt_2004_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054__entry__
      -- CP-element group 70: 	 branch_block_stmt_1739/merge_stmt_2018__exit__
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1739/if_stmt_2004_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1739/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1739/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1739/merge_stmt_2018_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1739/merge_stmt_2018_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1739/merge_stmt_2018_PhiAck/dummy
      -- 
    else_choice_transition_5100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2004_branch_ack_0, ack => convTransposeB_CP_4495_elements(70)); -- 
    rr_5116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(70), ack => type_cast_2032_inst_req_0); -- 
    cr_5135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(70), ack => type_cast_2048_inst_req_1); -- 
    cr_5121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(70), ack => type_cast_2032_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_sample_completed_
      -- 
    ra_5117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2032_inst_ack_0, ack => convTransposeB_CP_4495_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2032_update_completed_
      -- 
    ca_5122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2032_inst_ack_1, ack => convTransposeB_CP_4495_elements(72)); -- 
    rr_5130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(72), ack => type_cast_2048_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_sample_completed_
      -- 
    ra_5131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_0, ack => convTransposeB_CP_4495_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/$exit
      -- CP-element group 74: 	 branch_block_stmt_1739/R_cmp117_2056_place
      -- CP-element group 74: 	 branch_block_stmt_1739/if_stmt_2055__entry__
      -- CP-element group 74: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054__exit__
      -- CP-element group 74: 	 branch_block_stmt_1739/if_stmt_2055_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1739/if_stmt_2055_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1739/if_stmt_2055_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1739/if_stmt_2055_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1739/if_stmt_2055_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1739/if_stmt_2055_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1739/assign_stmt_2024_to_assign_stmt_2054/type_cast_2048_update_completed_
      -- 
    ca_5136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_1, ack => convTransposeB_CP_4495_elements(74)); -- 
    branch_req_5144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(74), ack => if_stmt_2055_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1739/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1739/merge_stmt_2089_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1739/assign_stmt_2094__entry__
      -- CP-element group 75: 	 branch_block_stmt_1739/merge_stmt_2089__exit__
      -- CP-element group 75: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1739/assign_stmt_2094/$entry
      -- CP-element group 75: 	 branch_block_stmt_1739/if_stmt_2055_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1739/if_stmt_2055_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1739/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1739/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1739/merge_stmt_2089_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1739/merge_stmt_2089_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1739/merge_stmt_2089_PhiAck/dummy
      -- 
    if_choice_transition_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2055_branch_ack_1, ack => convTransposeB_CP_4495_elements(75)); -- 
    req_5169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(75), ack => WPIPE_Block1_done_2091_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	111 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1739/if_stmt_2055_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1739/if_stmt_2055_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2062/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$entry
      -- 
    else_choice_transition_5153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2055_branch_ack_0, ack => convTransposeB_CP_4495_elements(76)); -- 
    rr_5371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(76), ack => type_cast_2080_inst_req_0); -- 
    cr_5376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(76), ack => type_cast_2080_inst_req_1); -- 
    rr_5394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(76), ack => type_cast_2074_inst_req_0); -- 
    cr_5399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(76), ack => type_cast_2074_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Update/req
      -- 
    ack_5170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2091_inst_ack_0, ack => convTransposeB_CP_4495_elements(77)); -- 
    req_5174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(77), ack => WPIPE_Block1_done_2091_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1739/merge_stmt_2096_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1739/assign_stmt_2094/$exit
      -- CP-element group 78: 	 branch_block_stmt_1739/merge_stmt_2096__exit__
      -- CP-element group 78: 	 branch_block_stmt_1739/return__
      -- CP-element group 78: 	 branch_block_stmt_1739/$exit
      -- CP-element group 78: 	 branch_block_stmt_1739/assign_stmt_2094__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1739/branch_block_stmt_1739__exit__
      -- CP-element group 78: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1739/assign_stmt_2094/WPIPE_Block1_done_2091_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1739/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1739/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1739/merge_stmt_2096_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1739/merge_stmt_2096_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1739/merge_stmt_2096_PhiAck/dummy
      -- 
    ack_5175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2091_inst_ack_1, ack => convTransposeB_CP_4495_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Sample/ra
      -- 
    ra_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1880_inst_ack_0, ack => convTransposeB_CP_4495_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/Update/ca
      -- 
    ca_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1880_inst_ack_1, ack => convTransposeB_CP_4495_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/$exit
      -- CP-element group 81: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/$exit
      -- CP-element group 81: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1880/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_req
      -- 
    phi_stmt_1875_req_5201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1875_req_5201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(81), ack => phi_stmt_1875_req_1); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(79) & convTransposeB_CP_4495_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1868/$exit
      -- CP-element group 82: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1872_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_req
      -- 
    phi_stmt_1868_req_5209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_req_5209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(82), ack => phi_stmt_1868_req_0); -- 
    -- Element group convTransposeB_CP_4495_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4495_elements(43), ack => convTransposeB_CP_4495_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1861/$exit
      -- CP-element group 83: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1865_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_req
      -- 
    phi_stmt_1861_req_5217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1861_req_5217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(83), ack => phi_stmt_1861_req_0); -- 
    -- Element group convTransposeB_CP_4495_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4495_elements(43), ack => convTransposeB_CP_4495_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1854/$exit
      -- CP-element group 84: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_req
      -- 
    phi_stmt_1854_req_5225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_req_5225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(84), ack => phi_stmt_1854_req_1); -- 
    -- Element group convTransposeB_CP_4495_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4495_elements(43), ack => convTransposeB_CP_4495_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1739/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(81) & convTransposeB_CP_4495_elements(82) & convTransposeB_CP_4495_elements(83) & convTransposeB_CP_4495_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Sample/ra
      -- 
    ra_5245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1878_inst_ack_0, ack => convTransposeB_CP_4495_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/Update/ca
      -- 
    ca_5250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1878_inst_ack_1, ack => convTransposeB_CP_4495_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/$exit
      -- CP-element group 88: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/$exit
      -- CP-element group 88: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1878/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_req
      -- 
    phi_stmt_1875_req_5251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1875_req_5251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(88), ack => phi_stmt_1875_req_0); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(86) & convTransposeB_CP_4495_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/ra
      -- 
    ra_5268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1874_inst_ack_0, ack => convTransposeB_CP_4495_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/ca
      -- 
    ca_5273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1874_inst_ack_1, ack => convTransposeB_CP_4495_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/$exit
      -- CP-element group 91: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/$exit
      -- CP-element group 91: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_req
      -- 
    phi_stmt_1868_req_5274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_req_5274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(91), ack => phi_stmt_1868_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(89) & convTransposeB_CP_4495_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Sample/ra
      -- 
    ra_5291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_0, ack => convTransposeB_CP_4495_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/Update/ca
      -- 
    ca_5296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_1, ack => convTransposeB_CP_4495_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/$exit
      -- CP-element group 94: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/$exit
      -- CP-element group 94: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_sources/type_cast_1867/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1861/phi_stmt_1861_req
      -- 
    phi_stmt_1861_req_5297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1861_req_5297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(94), ack => phi_stmt_1861_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(92) & convTransposeB_CP_4495_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/ra
      -- 
    ra_5314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_0, ack => convTransposeB_CP_4495_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/ca
      -- 
    ca_5319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_1, ack => convTransposeB_CP_4495_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/$exit
      -- CP-element group 97: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/$exit
      -- CP-element group 97: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1854/phi_stmt_1854_req
      -- 
    phi_stmt_1854_req_5320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_req_5320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(97), ack => phi_stmt_1854_req_0); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(95) & convTransposeB_CP_4495_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1739/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(88) & convTransposeB_CP_4495_elements(91) & convTransposeB_CP_4495_elements(94) & convTransposeB_CP_4495_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1739/merge_stmt_1853_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_1739/merge_stmt_1853_PhiAck/$entry
      -- 
    convTransposeB_CP_4495_elements(99) <= OrReduce(convTransposeB_CP_4495_elements(85) & convTransposeB_CP_4495_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1739/merge_stmt_1853_PhiAck/phi_stmt_1854_ack
      -- 
    phi_stmt_1854_ack_5325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1854_ack_0, ack => convTransposeB_CP_4495_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1739/merge_stmt_1853_PhiAck/phi_stmt_1861_ack
      -- 
    phi_stmt_1861_ack_5326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1861_ack_0, ack => convTransposeB_CP_4495_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1739/merge_stmt_1853_PhiAck/phi_stmt_1868_ack
      -- 
    phi_stmt_1868_ack_5327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1868_ack_0, ack => convTransposeB_CP_4495_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1739/merge_stmt_1853_PhiAck/phi_stmt_1875_ack
      -- 
    phi_stmt_1875_ack_5328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1875_ack_0, ack => convTransposeB_CP_4495_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003__entry__
      -- CP-element group 104: 	 branch_block_stmt_1739/merge_stmt_1853__exit__
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1983_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1991_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1964_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/ptr_deref_1986_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1959_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/array_obj_ref_1982_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1915_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1919_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1923_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/type_cast_1953_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1739/assign_stmt_1887_to_assign_stmt_2003/addr_of_1960_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/merge_stmt_1853_PhiAck/$exit
      -- 
    cr_5068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => ptr_deref_1986_store_0_req_1); -- 
    req_4922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => addr_of_1960_final_reg_req_1); -- 
    rr_5077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1991_inst_req_0); -- 
    req_5018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => addr_of_1983_final_reg_req_1); -- 
    cr_5082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1991_inst_req_1); -- 
    cr_4967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => ptr_deref_1964_load_0_req_1); -- 
    req_5003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => array_obj_ref_1982_index_offset_req_1); -- 
    req_4907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => array_obj_ref_1959_index_offset_req_1); -- 
    rr_4829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1915_inst_req_0); -- 
    cr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1915_inst_req_1); -- 
    rr_4843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1919_inst_req_0); -- 
    cr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1919_inst_req_1); -- 
    rr_4857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1923_inst_req_0); -- 
    cr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1923_inst_req_1); -- 
    rr_4871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1953_inst_req_0); -- 
    cr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(104), ack => type_cast_1953_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(100) & convTransposeB_CP_4495_elements(101) & convTransposeB_CP_4495_elements(102) & convTransposeB_CP_4495_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Sample/ra
      -- 
    ra_5372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2080_inst_ack_0, ack => convTransposeB_CP_4495_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/Update/ca
      -- 
    ca_5377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2080_inst_ack_1, ack => convTransposeB_CP_4495_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/$exit
      -- CP-element group 107: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/$exit
      -- CP-element group 107: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2080/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_req
      -- 
    phi_stmt_2075_req_5378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2075_req_5378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(107), ack => phi_stmt_2075_req_1); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(105) & convTransposeB_CP_4495_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Sample/ra
      -- 
    ra_5395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2074_inst_ack_0, ack => convTransposeB_CP_4495_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/Update/ca
      -- 
    ca_5400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2074_inst_ack_1, ack => convTransposeB_CP_4495_elements(109)); -- 
    -- CP-element group 110:  join  transition  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/$exit
      -- CP-element group 110: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/$exit
      -- CP-element group 110: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/$exit
      -- CP-element group 110: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2074/SplitProtocol/$exit
      -- CP-element group 110: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_req
      -- 
    phi_stmt_2069_req_5401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2069_req_5401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(110), ack => phi_stmt_2069_req_1); -- 
    convTransposeB_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(108) & convTransposeB_CP_4495_elements(109);
      gj_convTransposeB_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  output  delay-element  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	76 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2062/$exit
      -- CP-element group 111: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2068_konst_delay_trans
      -- CP-element group 111: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_req
      -- 
    phi_stmt_2062_req_5409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2062_req_5409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(111), ack => phi_stmt_2062_req_1); -- 
    -- Element group convTransposeB_CP_4495_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => convTransposeB_CP_4495_elements(76), ack => convTransposeB_CP_4495_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1739/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(107) & convTransposeB_CP_4495_elements(110) & convTransposeB_CP_4495_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Sample/ra
      -- 
    ra_5429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2078_inst_ack_0, ack => convTransposeB_CP_4495_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/Update/ca
      -- 
    ca_5434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2078_inst_ack_1, ack => convTransposeB_CP_4495_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/$exit
      -- CP-element group 115: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/$exit
      -- CP-element group 115: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_sources/type_cast_2078/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2075/phi_stmt_2075_req
      -- 
    phi_stmt_2075_req_5435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2075_req_5435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(115), ack => phi_stmt_2075_req_0); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(113) & convTransposeB_CP_4495_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Sample/ra
      -- 
    ra_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2072_inst_ack_0, ack => convTransposeB_CP_4495_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/Update/ca
      -- 
    ca_5457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2072_inst_ack_1, ack => convTransposeB_CP_4495_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/$exit
      -- CP-element group 118: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/$exit
      -- CP-element group 118: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_sources/type_cast_2072/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2069/phi_stmt_2069_req
      -- 
    phi_stmt_2069_req_5458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2069_req_5458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(118), ack => phi_stmt_2069_req_0); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(116) & convTransposeB_CP_4495_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/ra
      -- 
    ra_5475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_0, ack => convTransposeB_CP_4495_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/ca
      -- 
    ca_5480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_1, ack => convTransposeB_CP_4495_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/$exit
      -- CP-element group 121: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/$exit
      -- CP-element group 121: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2062/phi_stmt_2062_req
      -- 
    phi_stmt_2062_req_5481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2062_req_5481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4495_elements(121), ack => phi_stmt_2062_req_0); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(119) & convTransposeB_CP_4495_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1739/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(115) & convTransposeB_CP_4495_elements(118) & convTransposeB_CP_4495_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1739/merge_stmt_2061_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_1739/merge_stmt_2061_PhiAck/$entry
      -- 
    convTransposeB_CP_4495_elements(123) <= OrReduce(convTransposeB_CP_4495_elements(112) & convTransposeB_CP_4495_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1739/merge_stmt_2061_PhiAck/phi_stmt_2062_ack
      -- 
    phi_stmt_2062_ack_5486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2062_ack_0, ack => convTransposeB_CP_4495_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1739/merge_stmt_2061_PhiAck/phi_stmt_2069_ack
      -- 
    phi_stmt_2069_ack_5487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2069_ack_0, ack => convTransposeB_CP_4495_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1739/merge_stmt_2061_PhiAck/phi_stmt_2075_ack
      -- 
    phi_stmt_2075_ack_5488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2075_ack_0, ack => convTransposeB_CP_4495_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1739/merge_stmt_2061_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4495_elements(124) & convTransposeB_CP_4495_elements(125) & convTransposeB_CP_4495_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4495_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_1981_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_1981_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1958_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1958_scaled : std_logic_vector(13 downto 0);
    signal add45_1813 : std_logic_vector(15 downto 0);
    signal add58_1824 : std_logic_vector(15 downto 0);
    signal add77_1934 : std_logic_vector(63 downto 0);
    signal add79_1944 : std_logic_vector(63 downto 0);
    signal add91_1998 : std_logic_vector(31 downto 0);
    signal add98_2016 : std_logic_vector(15 downto 0);
    signal add_1791 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1892 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1959_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_1961 : std_logic_vector(31 downto 0);
    signal arrayidx87_1984 : std_logic_vector(31 downto 0);
    signal call11_1760 : std_logic_vector(15 downto 0);
    signal call13_1763 : std_logic_vector(15 downto 0);
    signal call14_1766 : std_logic_vector(15 downto 0);
    signal call15_1769 : std_logic_vector(15 downto 0);
    signal call16_1782 : std_logic_vector(15 downto 0);
    signal call18_1794 : std_logic_vector(15 downto 0);
    signal call1_1745 : std_logic_vector(15 downto 0);
    signal call20_1797 : std_logic_vector(15 downto 0);
    signal call22_1800 : std_logic_vector(15 downto 0);
    signal call3_1748 : std_logic_vector(15 downto 0);
    signal call5_1751 : std_logic_vector(15 downto 0);
    signal call7_1754 : std_logic_vector(15 downto 0);
    signal call9_1757 : std_logic_vector(15 downto 0);
    signal call_1742 : std_logic_vector(15 downto 0);
    signal cmp106_2029 : std_logic_vector(0 downto 0);
    signal cmp117_2054 : std_logic_vector(0 downto 0);
    signal cmp_2003 : std_logic_vector(0 downto 0);
    signal conv112_2049 : std_logic_vector(31 downto 0);
    signal conv115_1845 : std_logic_vector(31 downto 0);
    signal conv17_1786 : std_logic_vector(31 downto 0);
    signal conv65_1916 : std_logic_vector(63 downto 0);
    signal conv68_1833 : std_logic_vector(63 downto 0);
    signal conv70_1920 : std_logic_vector(63 downto 0);
    signal conv73_1837 : std_logic_vector(63 downto 0);
    signal conv75_1924 : std_logic_vector(63 downto 0);
    signal conv90_1992 : std_logic_vector(31 downto 0);
    signal conv94_1841 : std_logic_vector(31 downto 0);
    signal conv_1773 : std_logic_vector(31 downto 0);
    signal idxprom86_1977 : std_logic_vector(63 downto 0);
    signal idxprom_1954 : std_logic_vector(63 downto 0);
    signal inc110_2033 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2038 : std_logic_vector(15 downto 0);
    signal inc_2024 : std_logic_vector(15 downto 0);
    signal indvar_1854 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2087 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2075 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1875 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2069 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1868 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2045 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2062 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1861 : std_logic_vector(15 downto 0);
    signal mul54_1907 : std_logic_vector(15 downto 0);
    signal mul76_1929 : std_logic_vector(63 downto 0);
    signal mul78_1939 : std_logic_vector(63 downto 0);
    signal mul_1897 : std_logic_vector(15 downto 0);
    signal ptr_deref_1964_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1964_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1964_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1964_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1964_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1986_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1986_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1779 : std_logic_vector(31 downto 0);
    signal shr116132_1851 : std_logic_vector(31 downto 0);
    signal shr131_1807 : std_logic_vector(15 downto 0);
    signal shr81_1950 : std_logic_vector(31 downto 0);
    signal shr85_1971 : std_logic_vector(63 downto 0);
    signal sub48_1902 : std_logic_vector(15 downto 0);
    signal sub61_1829 : std_logic_vector(15 downto 0);
    signal sub62_1912 : std_logic_vector(15 downto 0);
    signal sub_1818 : std_logic_vector(15 downto 0);
    signal tmp1_1887 : std_logic_vector(31 downto 0);
    signal tmp83_1965 : std_logic_vector(63 downto 0);
    signal type_cast_1777_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1805_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1811_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1822_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1849_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1857_wire : std_logic_vector(31 downto 0);
    signal type_cast_1860_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1865_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1867_wire : std_logic_vector(15 downto 0);
    signal type_cast_1872_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1874_wire : std_logic_vector(15 downto 0);
    signal type_cast_1878_wire : std_logic_vector(15 downto 0);
    signal type_cast_1880_wire : std_logic_vector(15 downto 0);
    signal type_cast_1885_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1948_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1969_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1975_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1996_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2014_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2022_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2042_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2065_wire : std_logic_vector(15 downto 0);
    signal type_cast_2068_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2072_wire : std_logic_vector(15 downto 0);
    signal type_cast_2074_wire : std_logic_vector(15 downto 0);
    signal type_cast_2078_wire : std_logic_vector(15 downto 0);
    signal type_cast_2080_wire : std_logic_vector(15 downto 0);
    signal type_cast_2085_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2093_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1959_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1959_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1959_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1959_resized_base_address <= "00000000000000";
    array_obj_ref_1982_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1982_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1982_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1982_resized_base_address <= "00000000000000";
    ptr_deref_1964_word_offset_0 <= "00000000000000";
    ptr_deref_1986_word_offset_0 <= "00000000000000";
    type_cast_1777_wire_constant <= "00000000000000000000000000010000";
    type_cast_1805_wire_constant <= "0000000000000010";
    type_cast_1811_wire_constant <= "1111111111111111";
    type_cast_1822_wire_constant <= "1111111111111111";
    type_cast_1849_wire_constant <= "00000000000000000000000000000001";
    type_cast_1860_wire_constant <= "00000000000000000000000000000000";
    type_cast_1865_wire_constant <= "0000000000000000";
    type_cast_1872_wire_constant <= "0000000000000000";
    type_cast_1885_wire_constant <= "00000000000000000000000000000100";
    type_cast_1948_wire_constant <= "00000000000000000000000000000010";
    type_cast_1969_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1975_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1996_wire_constant <= "00000000000000000000000000000100";
    type_cast_2014_wire_constant <= "0000000000000100";
    type_cast_2022_wire_constant <= "0000000000000001";
    type_cast_2042_wire_constant <= "0000000000000000";
    type_cast_2068_wire_constant <= "0000000000000000";
    type_cast_2085_wire_constant <= "00000000000000000000000000000001";
    type_cast_2093_wire_constant <= "0000000000000001";
    phi_stmt_1854: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1857_wire & type_cast_1860_wire_constant;
      req <= phi_stmt_1854_req_0 & phi_stmt_1854_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1854",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1854_ack_0,
          idata => idata,
          odata => indvar_1854,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1854
    phi_stmt_1861: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1865_wire_constant & type_cast_1867_wire;
      req <= phi_stmt_1861_req_0 & phi_stmt_1861_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1861",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1861_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1861,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1861
    phi_stmt_1868: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1872_wire_constant & type_cast_1874_wire;
      req <= phi_stmt_1868_req_0 & phi_stmt_1868_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1868",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1868_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1868,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1868
    phi_stmt_1875: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1878_wire & type_cast_1880_wire;
      req <= phi_stmt_1875_req_0 & phi_stmt_1875_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1875",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1875_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1875,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1875
    phi_stmt_2062: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2065_wire & type_cast_2068_wire_constant;
      req <= phi_stmt_2062_req_0 & phi_stmt_2062_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2062",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2062_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2062,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2062
    phi_stmt_2069: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2072_wire & type_cast_2074_wire;
      req <= phi_stmt_2069_req_0 & phi_stmt_2069_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2069",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2069_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2069,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2069
    phi_stmt_2075: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2078_wire & type_cast_2080_wire;
      req <= phi_stmt_2075_req_0 & phi_stmt_2075_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2075",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2075_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2075,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2075
    -- flow-through select operator MUX_2044_inst
    input_dim1x_x2_2045 <= type_cast_2042_wire_constant when (cmp106_2029(0) /=  '0') else inc_2024;
    addr_of_1960_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1960_final_reg_req_0;
      addr_of_1960_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1960_final_reg_req_1;
      addr_of_1960_final_reg_ack_1<= rack(0);
      addr_of_1960_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1960_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1959_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1961,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1983_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1983_final_reg_req_0;
      addr_of_1983_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1983_final_reg_req_1;
      addr_of_1983_final_reg_ack_1<= rack(0);
      addr_of_1983_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1983_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1982_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_1984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1772_inst_req_0;
      type_cast_1772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1772_inst_req_1;
      type_cast_1772_inst_ack_1<= rack(0);
      type_cast_1772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1785_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1785_inst_req_0;
      type_cast_1785_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1785_inst_req_1;
      type_cast_1785_inst_ack_1<= rack(0);
      type_cast_1785_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1785_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1786,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1832_inst_req_0;
      type_cast_1832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1832_inst_req_1;
      type_cast_1832_inst_ack_1<= rack(0);
      type_cast_1832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1800,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1836_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1836_inst_req_0;
      type_cast_1836_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1836_inst_req_1;
      type_cast_1836_inst_ack_1<= rack(0);
      type_cast_1836_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1836_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1837,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1840_inst_req_0;
      type_cast_1840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1840_inst_req_1;
      type_cast_1840_inst_ack_1<= rack(0);
      type_cast_1840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1841,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1844_inst_req_0;
      type_cast_1844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1844_inst_req_1;
      type_cast_1844_inst_ack_1<= rack(0);
      type_cast_1844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1857_inst_req_0;
      type_cast_1857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1857_inst_req_1;
      type_cast_1857_inst_ack_1<= rack(0);
      type_cast_1857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2087,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1857_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1867_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1867_inst_req_0;
      type_cast_1867_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1867_inst_req_1;
      type_cast_1867_inst_ack_1<= rack(0);
      type_cast_1867_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1867_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2062,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1867_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1874_inst_req_0;
      type_cast_1874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1874_inst_req_1;
      type_cast_1874_inst_ack_1<= rack(0);
      type_cast_1874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2069,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1874_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1878_inst_req_0;
      type_cast_1878_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1878_inst_req_1;
      type_cast_1878_inst_ack_1<= rack(0);
      type_cast_1878_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1878_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2075,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1878_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1880_inst_req_0;
      type_cast_1880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1880_inst_req_1;
      type_cast_1880_inst_ack_1<= rack(0);
      type_cast_1880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1880_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1915_inst_req_0;
      type_cast_1915_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1915_inst_req_1;
      type_cast_1915_inst_ack_1<= rack(0);
      type_cast_1915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1915_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_1916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1919_inst_req_0;
      type_cast_1919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1919_inst_req_1;
      type_cast_1919_inst_ack_1<= rack(0);
      type_cast_1919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_1912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1920,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1923_inst_req_0;
      type_cast_1923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1923_inst_req_1;
      type_cast_1923_inst_ack_1<= rack(0);
      type_cast_1923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_1902,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1924,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1953_inst_req_0;
      type_cast_1953_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1953_inst_req_1;
      type_cast_1953_inst_ack_1<= rack(0);
      type_cast_1953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_1950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1991_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1991_inst_req_0;
      type_cast_1991_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1991_inst_req_1;
      type_cast_1991_inst_ack_1<= rack(0);
      type_cast_1991_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1991_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1992,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2032_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2032_inst_req_0;
      type_cast_2032_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2032_inst_req_1;
      type_cast_2032_inst_ack_1<= rack(0);
      type_cast_2032_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2032_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2033,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2048_inst_req_0;
      type_cast_2048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2048_inst_req_1;
      type_cast_2048_inst_ack_1<= rack(0);
      type_cast_2048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2038,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2065_inst_req_0;
      type_cast_2065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2065_inst_req_1;
      type_cast_2065_inst_ack_1<= rack(0);
      type_cast_2065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2016,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2065_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2072_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2072_inst_req_0;
      type_cast_2072_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2072_inst_req_1;
      type_cast_2072_inst_ack_1<= rack(0);
      type_cast_2072_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2072_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2072_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2074_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2074_inst_req_0;
      type_cast_2074_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2074_inst_req_1;
      type_cast_2074_inst_ack_1<= rack(0);
      type_cast_2074_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2074_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2074_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2078_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2078_inst_req_0;
      type_cast_2078_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2078_inst_req_1;
      type_cast_2078_inst_ack_1<= rack(0);
      type_cast_2078_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2078_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1875,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2078_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2080_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2080_inst_req_0;
      type_cast_2080_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2080_inst_req_1;
      type_cast_2080_inst_ack_1<= rack(0);
      type_cast_2080_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2080_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2038,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2080_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1959_index_1_rename
    process(R_idxprom_1958_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1958_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1958_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1959_index_1_resize
    process(idxprom_1954) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1954;
      ov := iv(13 downto 0);
      R_idxprom_1958_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1959_root_address_inst
    process(array_obj_ref_1959_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1959_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1959_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_index_1_rename
    process(R_idxprom86_1981_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_1981_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_1981_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_index_1_resize
    process(idxprom86_1977) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_1977;
      ov := iv(13 downto 0);
      R_idxprom86_1981_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_root_address_inst
    process(array_obj_ref_1982_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1982_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1982_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1964_addr_0
    process(ptr_deref_1964_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1964_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1964_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1964_base_resize
    process(arrayidx82_1961) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1961;
      ov := iv(13 downto 0);
      ptr_deref_1964_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1964_gather_scatter
    process(ptr_deref_1964_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1964_data_0;
      ov(63 downto 0) := iv;
      tmp83_1965 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1964_root_address_inst
    process(ptr_deref_1964_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1964_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1964_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_addr_0
    process(ptr_deref_1986_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1986_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1986_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_base_resize
    process(arrayidx87_1984) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_1984;
      ov := iv(13 downto 0);
      ptr_deref_1986_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_gather_scatter
    process(tmp83_1965) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_1965;
      ov(63 downto 0) := iv;
      ptr_deref_1986_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_root_address_inst
    process(ptr_deref_1986_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1986_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1986_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2004_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2003;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2004_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2004_branch_req_0,
          ack0 => if_stmt_2004_branch_ack_0,
          ack1 => if_stmt_2004_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2055_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2054;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2055_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2055_branch_req_0,
          ack0 => if_stmt_2055_branch_ack_0,
          ack1 => if_stmt_2055_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1812_inst
    process(call7_1754) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1754, type_cast_1811_wire_constant, tmp_var);
      add45_1813 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1823_inst
    process(call9_1757) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1757, type_cast_1822_wire_constant, tmp_var);
      add58_1824 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1901_inst
    process(sub_1818, mul_1897) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1818, mul_1897, tmp_var);
      sub48_1902 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1911_inst
    process(sub61_1829, mul54_1907) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1829, mul54_1907, tmp_var);
      sub62_1912 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2015_inst
    process(input_dim2x_x1_1861) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1861, type_cast_2014_wire_constant, tmp_var);
      add98_2016 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2023_inst
    process(input_dim1x_x1_1868) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1868, type_cast_2022_wire_constant, tmp_var);
      inc_2024 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2037_inst
    process(inc110_2033, input_dim0x_x2_1875) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2033, input_dim0x_x2_1875, tmp_var);
      inc110x_xinput_dim0x_x2_2038 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1891_inst
    process(add_1791, tmp1_1887) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1791, tmp1_1887, tmp_var);
      add_src_0x_x0_1892 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1997_inst
    process(conv90_1992) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_1992, type_cast_1996_wire_constant, tmp_var);
      add91_1998 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2086_inst
    process(indvar_1854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1854, type_cast_2085_wire_constant, tmp_var);
      indvarx_xnext_2087 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1933_inst
    process(mul76_1929, conv70_1920) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_1929, conv70_1920, tmp_var);
      add77_1934 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1943_inst
    process(mul78_1939, conv65_1916) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_1939, conv65_1916, tmp_var);
      add79_1944 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1976_inst
    process(shr85_1971) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_1971, type_cast_1975_wire_constant, tmp_var);
      idxprom86_1977 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2028_inst
    process(inc_2024, call1_1745) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2024, call1_1745, tmp_var);
      cmp106_2029 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2053_inst
    process(conv112_2049, shr116132_1851) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2049, shr116132_1851, tmp_var);
      cmp117_2054 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1806_inst
    process(call_1742) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1742, type_cast_1805_wire_constant, tmp_var);
      shr131_1807 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1850_inst
    process(conv115_1845) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1845, type_cast_1849_wire_constant, tmp_var);
      shr116132_1851 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1949_inst
    process(add_src_0x_x0_1892) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1892, type_cast_1948_wire_constant, tmp_var);
      shr81_1950 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1970_inst
    process(add79_1944) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_1944, type_cast_1969_wire_constant, tmp_var);
      shr85_1971 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1896_inst
    process(input_dim0x_x2_1875, call13_1763) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1875, call13_1763, tmp_var);
      mul_1897 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1906_inst
    process(input_dim1x_x1_1868, call13_1763) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1868, call13_1763, tmp_var);
      mul54_1907 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1886_inst
    process(indvar_1854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1854, type_cast_1885_wire_constant, tmp_var);
      tmp1_1887 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1928_inst
    process(conv75_1924, conv73_1837) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_1924, conv73_1837, tmp_var);
      mul76_1929 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1938_inst
    process(add77_1934, conv68_1833) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_1934, conv68_1833, tmp_var);
      mul78_1939 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1790_inst
    process(shl_1779, conv17_1786) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1779, conv17_1786, tmp_var);
      add_1791 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1778_inst
    process(conv_1773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1773, type_cast_1777_wire_constant, tmp_var);
      shl_1779 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1817_inst
    process(add45_1813, call14_1766) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1813, call14_1766, tmp_var);
      sub_1818 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1828_inst
    process(add58_1824, call14_1766) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1824, call14_1766, tmp_var);
      sub61_1829 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2002_inst
    process(add91_1998, conv94_1841) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_1998, conv94_1841, tmp_var);
      cmp_2003 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_1959_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1958_scaled;
      array_obj_ref_1959_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1959_index_offset_req_0;
      array_obj_ref_1959_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1959_index_offset_req_1;
      array_obj_ref_1959_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_1982_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_1981_scaled;
      array_obj_ref_1982_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1982_index_offset_req_0;
      array_obj_ref_1982_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1982_index_offset_req_1;
      array_obj_ref_1982_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_1964_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1964_load_0_req_0;
      ptr_deref_1964_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1964_load_0_req_1;
      ptr_deref_1964_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1964_word_address_0;
      ptr_deref_1964_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1986_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1986_store_0_req_0;
      ptr_deref_1986_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1986_store_0_req_1;
      ptr_deref_1986_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1986_word_address_0;
      data_in <= ptr_deref_1986_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1741_inst RPIPE_Block1_start_1744_inst RPIPE_Block1_start_1747_inst RPIPE_Block1_start_1750_inst RPIPE_Block1_start_1753_inst RPIPE_Block1_start_1756_inst RPIPE_Block1_start_1759_inst RPIPE_Block1_start_1762_inst RPIPE_Block1_start_1765_inst RPIPE_Block1_start_1768_inst RPIPE_Block1_start_1781_inst RPIPE_Block1_start_1793_inst RPIPE_Block1_start_1796_inst RPIPE_Block1_start_1799_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1741_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1744_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1747_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1750_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1753_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1756_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1759_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1762_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1765_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1768_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1781_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1793_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1796_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1799_inst_req_0;
      RPIPE_Block1_start_1741_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1744_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1747_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1750_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1753_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1756_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1759_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1762_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1765_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1768_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1781_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1793_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1796_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1799_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1741_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1744_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1747_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1750_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1753_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1756_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1759_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1762_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1765_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1768_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1781_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1793_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1796_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1799_inst_req_1;
      RPIPE_Block1_start_1741_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1744_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1747_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1750_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1753_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1756_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1759_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1762_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1765_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1768_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1781_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1793_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1796_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1799_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_1742 <= data_out(223 downto 208);
      call1_1745 <= data_out(207 downto 192);
      call3_1748 <= data_out(191 downto 176);
      call5_1751 <= data_out(175 downto 160);
      call7_1754 <= data_out(159 downto 144);
      call9_1757 <= data_out(143 downto 128);
      call11_1760 <= data_out(127 downto 112);
      call13_1763 <= data_out(111 downto 96);
      call14_1766 <= data_out(95 downto 80);
      call15_1769 <= data_out(79 downto 64);
      call16_1782 <= data_out(63 downto 48);
      call18_1794 <= data_out(47 downto 32);
      call20_1797 <= data_out(31 downto 16);
      call22_1800 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2091_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2091_inst_req_0;
      WPIPE_Block1_done_2091_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2091_inst_req_1;
      WPIPE_Block1_done_2091_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2093_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5505_start: Boolean;
  signal convTransposeC_CP_5505_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2420_inst_req_0 : boolean;
  signal ptr_deref_2358_store_0_req_1 : boolean;
  signal type_cast_2246_inst_ack_0 : boolean;
  signal type_cast_2404_inst_ack_1 : boolean;
  signal type_cast_2404_inst_req_1 : boolean;
  signal type_cast_2404_inst_ack_0 : boolean;
  signal type_cast_2404_inst_req_0 : boolean;
  signal type_cast_2239_inst_ack_0 : boolean;
  signal type_cast_2420_inst_ack_0 : boolean;
  signal phi_stmt_2233_req_0 : boolean;
  signal type_cast_2239_inst_req_0 : boolean;
  signal ptr_deref_2358_store_0_ack_0 : boolean;
  signal RPIPE_Block2_start_2108_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2108_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2108_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2108_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2105_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2105_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2105_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2105_inst_req_0 : boolean;
  signal addr_of_2355_final_reg_ack_0 : boolean;
  signal type_cast_2232_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2111_inst_ack_1 : boolean;
  signal type_cast_2232_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2111_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2111_inst_req_0 : boolean;
  signal addr_of_2355_final_reg_req_0 : boolean;
  signal phi_stmt_2247_req_1 : boolean;
  signal RPIPE_Block2_start_2102_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2102_inst_req_1 : boolean;
  signal type_cast_2232_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2102_inst_ack_0 : boolean;
  signal ptr_deref_2358_store_0_req_0 : boolean;
  signal RPIPE_Block2_start_2102_inst_req_0 : boolean;
  signal type_cast_2246_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2111_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2114_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2114_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2117_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2117_inst_ack_0 : boolean;
  signal type_cast_2252_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2114_inst_ack_0 : boolean;
  signal type_cast_2420_inst_req_1 : boolean;
  signal type_cast_2232_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2114_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2117_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2117_inst_req_1 : boolean;
  signal type_cast_2252_inst_ack_1 : boolean;
  signal type_cast_2246_inst_req_1 : boolean;
  signal phi_stmt_2226_req_1 : boolean;
  signal type_cast_2420_inst_ack_1 : boolean;
  signal phi_stmt_2226_req_0 : boolean;
  signal RPIPE_Block2_start_2120_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2120_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2120_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2463_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2120_inst_ack_1 : boolean;
  signal if_stmt_2376_branch_ack_0 : boolean;
  signal RPIPE_Block2_start_2123_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2463_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2123_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2123_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2123_inst_ack_1 : boolean;
  signal phi_stmt_2247_req_0 : boolean;
  signal RPIPE_Block2_start_2126_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2126_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2126_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2463_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2126_inst_ack_1 : boolean;
  signal type_cast_2250_inst_ack_1 : boolean;
  signal type_cast_2250_inst_req_1 : boolean;
  signal if_stmt_2376_branch_ack_1 : boolean;
  signal type_cast_2252_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2129_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2463_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2129_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2129_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2129_inst_ack_1 : boolean;
  signal type_cast_2250_inst_ack_0 : boolean;
  signal type_cast_2250_inst_req_0 : boolean;
  signal type_cast_2252_inst_req_0 : boolean;
  signal if_stmt_2376_branch_req_0 : boolean;
  signal type_cast_2133_inst_req_0 : boolean;
  signal type_cast_2133_inst_ack_0 : boolean;
  signal type_cast_2133_inst_req_1 : boolean;
  signal type_cast_2133_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2142_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2142_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2142_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2142_inst_ack_1 : boolean;
  signal array_obj_ref_2354_index_offset_ack_1 : boolean;
  signal array_obj_ref_2354_index_offset_req_1 : boolean;
  signal type_cast_2146_inst_req_0 : boolean;
  signal type_cast_2146_inst_ack_0 : boolean;
  signal type_cast_2146_inst_req_1 : boolean;
  signal type_cast_2146_inst_ack_1 : boolean;
  signal phi_stmt_2226_ack_0 : boolean;
  signal RPIPE_Block2_start_2154_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2154_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2154_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2154_inst_ack_1 : boolean;
  signal array_obj_ref_2354_index_offset_ack_0 : boolean;
  signal array_obj_ref_2354_index_offset_req_0 : boolean;
  signal RPIPE_Block2_start_2157_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2157_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2157_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2157_inst_ack_1 : boolean;
  signal type_cast_2363_inst_ack_1 : boolean;
  signal type_cast_2363_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2160_inst_req_0 : boolean;
  signal if_stmt_2427_branch_ack_0 : boolean;
  signal RPIPE_Block2_start_2160_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2160_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2160_inst_ack_1 : boolean;
  signal phi_stmt_2240_req_1 : boolean;
  signal type_cast_2246_inst_ack_1 : boolean;
  signal type_cast_2363_inst_ack_0 : boolean;
  signal type_cast_2193_inst_req_0 : boolean;
  signal if_stmt_2427_branch_ack_1 : boolean;
  signal type_cast_2193_inst_ack_0 : boolean;
  signal type_cast_2193_inst_req_1 : boolean;
  signal type_cast_2193_inst_ack_1 : boolean;
  signal type_cast_2363_inst_req_0 : boolean;
  signal type_cast_2197_inst_req_0 : boolean;
  signal type_cast_2197_inst_ack_0 : boolean;
  signal type_cast_2197_inst_req_1 : boolean;
  signal if_stmt_2427_branch_req_0 : boolean;
  signal type_cast_2197_inst_ack_1 : boolean;
  signal type_cast_2201_inst_req_0 : boolean;
  signal type_cast_2201_inst_ack_0 : boolean;
  signal phi_stmt_2233_req_1 : boolean;
  signal type_cast_2201_inst_req_1 : boolean;
  signal type_cast_2201_inst_ack_1 : boolean;
  signal ptr_deref_2358_store_0_ack_1 : boolean;
  signal type_cast_2239_inst_ack_1 : boolean;
  signal type_cast_2205_inst_req_0 : boolean;
  signal type_cast_2205_inst_ack_0 : boolean;
  signal type_cast_2239_inst_req_1 : boolean;
  signal type_cast_2205_inst_req_1 : boolean;
  signal type_cast_2205_inst_ack_1 : boolean;
  signal addr_of_2355_final_reg_ack_1 : boolean;
  signal phi_stmt_2240_req_0 : boolean;
  signal addr_of_2355_final_reg_req_1 : boolean;
  signal type_cast_2287_inst_req_0 : boolean;
  signal type_cast_2287_inst_ack_0 : boolean;
  signal type_cast_2287_inst_req_1 : boolean;
  signal type_cast_2287_inst_ack_1 : boolean;
  signal type_cast_2291_inst_req_0 : boolean;
  signal type_cast_2291_inst_ack_0 : boolean;
  signal type_cast_2291_inst_req_1 : boolean;
  signal type_cast_2291_inst_ack_1 : boolean;
  signal type_cast_2295_inst_req_0 : boolean;
  signal type_cast_2295_inst_ack_0 : boolean;
  signal type_cast_2295_inst_req_1 : boolean;
  signal type_cast_2295_inst_ack_1 : boolean;
  signal type_cast_2325_inst_req_0 : boolean;
  signal type_cast_2325_inst_ack_0 : boolean;
  signal type_cast_2325_inst_req_1 : boolean;
  signal type_cast_2325_inst_ack_1 : boolean;
  signal array_obj_ref_2331_index_offset_req_0 : boolean;
  signal array_obj_ref_2331_index_offset_ack_0 : boolean;
  signal array_obj_ref_2331_index_offset_req_1 : boolean;
  signal array_obj_ref_2331_index_offset_ack_1 : boolean;
  signal addr_of_2332_final_reg_req_0 : boolean;
  signal addr_of_2332_final_reg_ack_0 : boolean;
  signal addr_of_2332_final_reg_req_1 : boolean;
  signal addr_of_2332_final_reg_ack_1 : boolean;
  signal ptr_deref_2336_load_0_req_0 : boolean;
  signal ptr_deref_2336_load_0_ack_0 : boolean;
  signal ptr_deref_2336_load_0_req_1 : boolean;
  signal ptr_deref_2336_load_0_ack_1 : boolean;
  signal phi_stmt_2233_ack_0 : boolean;
  signal phi_stmt_2240_ack_0 : boolean;
  signal phi_stmt_2247_ack_0 : boolean;
  signal phi_stmt_2434_req_1 : boolean;
  signal type_cast_2444_inst_req_0 : boolean;
  signal type_cast_2444_inst_ack_0 : boolean;
  signal type_cast_2444_inst_req_1 : boolean;
  signal type_cast_2444_inst_ack_1 : boolean;
  signal phi_stmt_2441_req_0 : boolean;
  signal type_cast_2450_inst_req_0 : boolean;
  signal type_cast_2450_inst_ack_0 : boolean;
  signal type_cast_2450_inst_req_1 : boolean;
  signal type_cast_2450_inst_ack_1 : boolean;
  signal phi_stmt_2447_req_0 : boolean;
  signal type_cast_2437_inst_req_0 : boolean;
  signal type_cast_2437_inst_ack_0 : boolean;
  signal type_cast_2437_inst_req_1 : boolean;
  signal type_cast_2437_inst_ack_1 : boolean;
  signal phi_stmt_2434_req_0 : boolean;
  signal type_cast_2446_inst_req_0 : boolean;
  signal type_cast_2446_inst_ack_0 : boolean;
  signal type_cast_2446_inst_req_1 : boolean;
  signal type_cast_2446_inst_ack_1 : boolean;
  signal phi_stmt_2441_req_1 : boolean;
  signal type_cast_2452_inst_req_0 : boolean;
  signal type_cast_2452_inst_ack_0 : boolean;
  signal type_cast_2452_inst_req_1 : boolean;
  signal type_cast_2452_inst_ack_1 : boolean;
  signal phi_stmt_2447_req_1 : boolean;
  signal phi_stmt_2434_ack_0 : boolean;
  signal phi_stmt_2441_ack_0 : boolean;
  signal phi_stmt_2447_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5505_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5505_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5505_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5505_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5505: Block -- control-path 
    signal convTransposeC_CP_5505_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5505_elements(0) <= convTransposeC_CP_5505_start;
    convTransposeC_CP_5505_symbol <= convTransposeC_CP_5505_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161__entry__
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2100/branch_block_stmt_2100__entry__
      -- CP-element group 0: 	 branch_block_stmt_2100/$entry
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/$entry
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Update/cr
      -- 
    rr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(0), ack => RPIPE_Block2_start_2102_inst_req_0); -- 
    cr_5698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(0), ack => type_cast_2133_inst_req_1); -- 
    cr_5726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(0), ack => type_cast_2146_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2100/assign_stmt_2459__exit__
      -- CP-element group 1: 	 branch_block_stmt_2100/assign_stmt_2459__entry__
      -- CP-element group 1: 	 branch_block_stmt_2100/merge_stmt_2433__exit__
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/assign_stmt_2459/$exit
      -- CP-element group 1: 	 branch_block_stmt_2100/assign_stmt_2459/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/$entry
      -- 
    rr_6254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2239_inst_req_0); -- 
    cr_6328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2232_inst_req_1); -- 
    rr_6277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2246_inst_req_0); -- 
    rr_6323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2232_inst_req_0); -- 
    cr_6282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2246_inst_req_1); -- 
    cr_6305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2250_inst_req_1); -- 
    rr_6300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2250_inst_req_0); -- 
    cr_6259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(1), ack => type_cast_2239_inst_req_1); -- 
    convTransposeC_CP_5505_elements(1) <= convTransposeC_CP_5505_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_sample_completed_
      -- 
    ra_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2102_inst_ack_0, ack => convTransposeC_CP_5505_elements(2)); -- 
    cr_5558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(2), ack => RPIPE_Block2_start_2102_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2102_update_completed_
      -- 
    ca_5559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2102_inst_ack_1, ack => convTransposeC_CP_5505_elements(3)); -- 
    rr_5567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(3), ack => RPIPE_Block2_start_2105_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_sample_completed_
      -- 
    ra_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2105_inst_ack_0, ack => convTransposeC_CP_5505_elements(4)); -- 
    cr_5572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(4), ack => RPIPE_Block2_start_2105_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2105_update_completed_
      -- 
    ca_5573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2105_inst_ack_1, ack => convTransposeC_CP_5505_elements(5)); -- 
    rr_5581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(5), ack => RPIPE_Block2_start_2108_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_sample_completed_
      -- 
    ra_5582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2108_inst_ack_0, ack => convTransposeC_CP_5505_elements(6)); -- 
    cr_5586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(6), ack => RPIPE_Block2_start_2108_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2108_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_sample_start_
      -- 
    ca_5587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2108_inst_ack_1, ack => convTransposeC_CP_5505_elements(7)); -- 
    rr_5595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(7), ack => RPIPE_Block2_start_2111_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Sample/ra
      -- 
    ra_5596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2111_inst_ack_0, ack => convTransposeC_CP_5505_elements(8)); -- 
    cr_5600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(8), ack => RPIPE_Block2_start_2111_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2111_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Sample/$entry
      -- 
    ca_5601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2111_inst_ack_1, ack => convTransposeC_CP_5505_elements(9)); -- 
    rr_5609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(9), ack => RPIPE_Block2_start_2114_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Sample/ra
      -- 
    ra_5610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2114_inst_ack_0, ack => convTransposeC_CP_5505_elements(10)); -- 
    cr_5614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(10), ack => RPIPE_Block2_start_2114_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2114_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Sample/$entry
      -- 
    ca_5615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2114_inst_ack_1, ack => convTransposeC_CP_5505_elements(11)); -- 
    rr_5623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(11), ack => RPIPE_Block2_start_2117_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Update/cr
      -- 
    ra_5624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2117_inst_ack_0, ack => convTransposeC_CP_5505_elements(12)); -- 
    cr_5628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(12), ack => RPIPE_Block2_start_2117_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2117_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Sample/rr
      -- 
    ca_5629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2117_inst_ack_1, ack => convTransposeC_CP_5505_elements(13)); -- 
    rr_5637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(13), ack => RPIPE_Block2_start_2120_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Update/cr
      -- 
    ra_5638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2120_inst_ack_0, ack => convTransposeC_CP_5505_elements(14)); -- 
    cr_5642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(14), ack => RPIPE_Block2_start_2120_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2120_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Sample/rr
      -- 
    ca_5643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2120_inst_ack_1, ack => convTransposeC_CP_5505_elements(15)); -- 
    rr_5651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(15), ack => RPIPE_Block2_start_2123_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Update/cr
      -- 
    ra_5652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2123_inst_ack_0, ack => convTransposeC_CP_5505_elements(16)); -- 
    cr_5656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(16), ack => RPIPE_Block2_start_2123_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2123_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Sample/rr
      -- 
    ca_5657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2123_inst_ack_1, ack => convTransposeC_CP_5505_elements(17)); -- 
    rr_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(17), ack => RPIPE_Block2_start_2126_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Update/cr
      -- 
    ra_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2126_inst_ack_0, ack => convTransposeC_CP_5505_elements(18)); -- 
    cr_5670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(18), ack => RPIPE_Block2_start_2126_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2126_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Sample/rr
      -- 
    ca_5671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2126_inst_ack_1, ack => convTransposeC_CP_5505_elements(19)); -- 
    rr_5679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(19), ack => RPIPE_Block2_start_2129_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Update/cr
      -- 
    ra_5680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2129_inst_ack_0, ack => convTransposeC_CP_5505_elements(20)); -- 
    cr_5684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(20), ack => RPIPE_Block2_start_2129_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2129_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Sample/rr
      -- 
    ca_5685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2129_inst_ack_1, ack => convTransposeC_CP_5505_elements(21)); -- 
    rr_5693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(21), ack => type_cast_2133_inst_req_0); -- 
    rr_5707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(21), ack => RPIPE_Block2_start_2142_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Sample/ra
      -- 
    ra_5694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_0, ack => convTransposeC_CP_5505_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2133_Update/ca
      -- 
    ca_5699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_1, ack => convTransposeC_CP_5505_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Update/cr
      -- 
    ra_5708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2142_inst_ack_0, ack => convTransposeC_CP_5505_elements(24)); -- 
    cr_5712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(24), ack => RPIPE_Block2_start_2142_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2142_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Sample/rr
      -- 
    ca_5713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2142_inst_ack_1, ack => convTransposeC_CP_5505_elements(25)); -- 
    rr_5721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(25), ack => type_cast_2146_inst_req_0); -- 
    rr_5735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(25), ack => RPIPE_Block2_start_2154_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Sample/ra
      -- 
    ra_5722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_0, ack => convTransposeC_CP_5505_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/type_cast_2146_Update/ca
      -- 
    ca_5727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_1, ack => convTransposeC_CP_5505_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Update/cr
      -- 
    ra_5736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2154_inst_ack_0, ack => convTransposeC_CP_5505_elements(28)); -- 
    cr_5740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(28), ack => RPIPE_Block2_start_2154_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2154_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Sample/rr
      -- 
    ca_5741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2154_inst_ack_1, ack => convTransposeC_CP_5505_elements(29)); -- 
    rr_5749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(29), ack => RPIPE_Block2_start_2157_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Update/cr
      -- 
    ra_5750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2157_inst_ack_0, ack => convTransposeC_CP_5505_elements(30)); -- 
    cr_5754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(30), ack => RPIPE_Block2_start_2157_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2157_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Sample/rr
      -- 
    ca_5755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2157_inst_ack_1, ack => convTransposeC_CP_5505_elements(31)); -- 
    rr_5763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(31), ack => RPIPE_Block2_start_2160_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Update/cr
      -- 
    ra_5764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2160_inst_ack_0, ack => convTransposeC_CP_5505_elements(32)); -- 
    cr_5768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(32), ack => RPIPE_Block2_start_2160_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/RPIPE_Block2_start_2160_Update/ca
      -- 
    ca_5769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2160_inst_ack_1, ack => convTransposeC_CP_5505_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223__entry__
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161__exit__
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2103_to_assign_stmt_2161/$exit
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Update/cr
      -- 
    rr_5780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2193_inst_req_0); -- 
    cr_5785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2193_inst_req_1); -- 
    rr_5794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2197_inst_req_0); -- 
    cr_5799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2197_inst_req_1); -- 
    rr_5808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2201_inst_req_0); -- 
    cr_5813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2201_inst_req_1); -- 
    rr_5822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2205_inst_req_0); -- 
    cr_5827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(34), ack => type_cast_2205_inst_req_1); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(23) & convTransposeC_CP_5505_elements(27) & convTransposeC_CP_5505_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Sample/ra
      -- 
    ra_5781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_0, ack => convTransposeC_CP_5505_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2193_Update/ca
      -- 
    ca_5786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_1, ack => convTransposeC_CP_5505_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Sample/ra
      -- 
    ra_5795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_0, ack => convTransposeC_CP_5505_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2197_Update/ca
      -- 
    ca_5800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_1, ack => convTransposeC_CP_5505_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Sample/ra
      -- 
    ra_5809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2201_inst_ack_0, ack => convTransposeC_CP_5505_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2201_Update/ca
      -- 
    ca_5814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2201_inst_ack_1, ack => convTransposeC_CP_5505_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Sample/ra
      -- 
    ra_5823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2205_inst_ack_0, ack => convTransposeC_CP_5505_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/type_cast_2205_Update/ca
      -- 
    ca_5828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2205_inst_ack_1, ack => convTransposeC_CP_5505_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2226/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223__exit__
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2233/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/assign_stmt_2168_to_assign_stmt_2223/$exit
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/$entry
      -- 
    cr_6225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(43), ack => type_cast_2252_inst_req_1); -- 
    rr_6220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(43), ack => type_cast_2252_inst_req_0); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(36) & convTransposeC_CP_5505_elements(38) & convTransposeC_CP_5505_elements(40) & convTransposeC_CP_5505_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Sample/ra
      -- 
    ra_5840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_0, ack => convTransposeC_CP_5505_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Update/ca
      -- 
    ca_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_1, ack => convTransposeC_CP_5505_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Sample/ra
      -- 
    ra_5854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2291_inst_ack_0, ack => convTransposeC_CP_5505_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Update/ca
      -- 
    ca_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2291_inst_ack_1, ack => convTransposeC_CP_5505_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Sample/ra
      -- 
    ra_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_0, ack => convTransposeC_CP_5505_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Update/ca
      -- 
    ca_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_1, ack => convTransposeC_CP_5505_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Sample/ra
      -- 
    ra_5882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2325_inst_ack_0, ack => convTransposeC_CP_5505_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Sample/req
      -- 
    ca_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2325_inst_ack_1, ack => convTransposeC_CP_5505_elements(51)); -- 
    req_5912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(51), ack => array_obj_ref_2331_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Sample/ack
      -- 
    ack_5913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2331_index_offset_ack_0, ack => convTransposeC_CP_5505_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_request/req
      -- 
    ack_5918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2331_index_offset_ack_1, ack => convTransposeC_CP_5505_elements(53)); -- 
    req_5927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(53), ack => addr_of_2332_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_request/ack
      -- 
    ack_5928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2332_final_reg_ack_0, ack => convTransposeC_CP_5505_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/word_access_start/word_0/rr
      -- 
    ack_5933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2332_final_reg_ack_1, ack => convTransposeC_CP_5505_elements(55)); -- 
    rr_5966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(55), ack => ptr_deref_2336_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Sample/word_access_start/word_0/ra
      -- 
    ra_5967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2336_load_0_ack_0, ack => convTransposeC_CP_5505_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/ptr_deref_2336_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/ptr_deref_2336_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/ptr_deref_2336_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/ptr_deref_2336_Merge/merge_ack
      -- 
    ca_5978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2336_load_0_ack_1, ack => convTransposeC_CP_5505_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_index_resize_1/index_resize_ack
      -- 
    req_6008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(58), ack => array_obj_ref_2354_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(45) & convTransposeC_CP_5505_elements(47) & convTransposeC_CP_5505_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Sample/$exit
      -- 
    ack_6009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2354_index_offset_ack_0, ack => convTransposeC_CP_5505_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_request/req
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_offset_calculated
      -- 
    ack_6014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2354_index_offset_ack_1, ack => convTransposeC_CP_5505_elements(60)); -- 
    req_6023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(60), ack => addr_of_2355_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_request/ack
      -- CP-element group 61: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_sample_completed_
      -- 
    ack_6024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2355_final_reg_ack_0, ack => convTransposeC_CP_5505_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_update_completed_
      -- 
    ack_6029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2355_final_reg_ack_1, ack => convTransposeC_CP_5505_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/ptr_deref_2358_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/ptr_deref_2358_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/ptr_deref_2358_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/ptr_deref_2358_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/word_access_start/word_0/rr
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_sample_start_
      -- 
    rr_6067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(63), ack => ptr_deref_2358_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(57) & convTransposeC_CP_5505_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/word_access_start/word_0/ra
      -- CP-element group 64: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_sample_completed_
      -- 
    ra_6068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2358_store_0_ack_0, ack => convTransposeC_CP_5505_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/word_access_complete/word_0/ca
      -- 
    ca_6079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2358_store_0_ack_1, ack => convTransposeC_CP_5505_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_sample_completed_
      -- 
    ra_6088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_0, ack => convTransposeC_CP_5505_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_update_completed_
      -- 
    ca_6093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_1, ack => convTransposeC_CP_5505_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2100/if_stmt_2376__entry__
      -- CP-element group 68: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375__exit__
      -- CP-element group 68: 	 branch_block_stmt_2100/if_stmt_2376_else_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2100/if_stmt_2376_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2100/if_stmt_2376_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2100/if_stmt_2376_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2100/if_stmt_2376_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2100/if_stmt_2376_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2100/R_cmp_2377_place
      -- CP-element group 68: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/$exit
      -- 
    branch_req_6101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(68), ack => if_stmt_2376_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(52) & convTransposeC_CP_5505_elements(59) & convTransposeC_CP_5505_elements(65) & convTransposeC_CP_5505_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2100/merge_stmt_2382__exit__
      -- CP-element group 69: 	 branch_block_stmt_2100/merge_stmt_2382_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2100/assign_stmt_2388/$exit
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2100/assign_stmt_2388__exit__
      -- CP-element group 69: 	 branch_block_stmt_2100/assign_stmt_2388__entry__
      -- CP-element group 69: 	 branch_block_stmt_2100/assign_stmt_2388/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/if_stmt_2376_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2100/if_stmt_2376_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2100/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2100/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2100/merge_stmt_2382_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/merge_stmt_2382_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2100/merge_stmt_2382_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2376_branch_ack_1, ack => convTransposeC_CP_5505_elements(69)); -- 
    rr_6438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(69), ack => type_cast_2437_inst_req_0); -- 
    cr_6443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(69), ack => type_cast_2437_inst_req_1); -- 
    rr_6461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(69), ack => type_cast_2446_inst_req_0); -- 
    cr_6466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(69), ack => type_cast_2446_inst_req_1); -- 
    rr_6484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(69), ack => type_cast_2452_inst_req_0); -- 
    cr_6489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(69), ack => type_cast_2452_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/$entry
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2100/merge_stmt_2390_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426__entry__
      -- CP-element group 70: 	 branch_block_stmt_2100/merge_stmt_2390__exit__
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2100/if_stmt_2376_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2100/if_stmt_2376_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2100/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2100/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2100/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2100/merge_stmt_2390_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2100/merge_stmt_2390_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2100/merge_stmt_2390_PhiAck/dummy
      -- 
    else_choice_transition_6110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2376_branch_ack_0, ack => convTransposeC_CP_5505_elements(70)); -- 
    cr_6131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(70), ack => type_cast_2404_inst_req_1); -- 
    rr_6126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(70), ack => type_cast_2404_inst_req_0); -- 
    cr_6145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(70), ack => type_cast_2420_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_sample_completed_
      -- 
    ra_6127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_0, ack => convTransposeC_CP_5505_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2404_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Sample/$entry
      -- 
    ca_6132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_1, ack => convTransposeC_CP_5505_elements(72)); -- 
    rr_6140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(72), ack => type_cast_2420_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Sample/$exit
      -- 
    ra_6141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2420_inst_ack_0, ack => convTransposeC_CP_5505_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/$exit
      -- CP-element group 74: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2100/if_stmt_2427__entry__
      -- CP-element group 74: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426__exit__
      -- CP-element group 74: 	 branch_block_stmt_2100/if_stmt_2427_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2100/assign_stmt_2396_to_assign_stmt_2426/type_cast_2420_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2100/if_stmt_2427_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2100/R_cmp122_2428_place
      -- CP-element group 74: 	 branch_block_stmt_2100/if_stmt_2427_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2100/if_stmt_2427_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2100/if_stmt_2427_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2100/if_stmt_2427_eval_test/$entry
      -- 
    ca_6146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2420_inst_ack_1, ack => convTransposeC_CP_5505_elements(74)); -- 
    branch_req_6154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(74), ack => if_stmt_2427_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2100/merge_stmt_2461_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2100/assign_stmt_2466__entry__
      -- CP-element group 75: 	 branch_block_stmt_2100/merge_stmt_2461__exit__
      -- CP-element group 75: 	 branch_block_stmt_2100/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2100/assign_stmt_2466/$entry
      -- CP-element group 75: 	 branch_block_stmt_2100/if_stmt_2427_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2100/if_stmt_2427_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2100/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2100/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2100/merge_stmt_2461_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2100/merge_stmt_2461_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2100/merge_stmt_2461_PhiAck/dummy
      -- 
    if_choice_transition_6159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2427_branch_ack_1, ack => convTransposeC_CP_5505_elements(75)); -- 
    req_6179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(75), ack => WPIPE_Block2_done_2463_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2100/if_stmt_2427_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2100/if_stmt_2427_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2434/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2427_branch_ack_0, ack => convTransposeC_CP_5505_elements(76)); -- 
    rr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(76), ack => type_cast_2444_inst_req_0); -- 
    cr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(76), ack => type_cast_2444_inst_req_1); -- 
    rr_6412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(76), ack => type_cast_2450_inst_req_0); -- 
    cr_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(76), ack => type_cast_2450_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Update/req
      -- CP-element group 77: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_sample_completed_
      -- 
    ack_6180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2463_inst_ack_0, ack => convTransposeC_CP_5505_elements(77)); -- 
    req_6184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(77), ack => WPIPE_Block2_done_2463_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_2100/merge_stmt_2468__exit__
      -- CP-element group 78: 	 branch_block_stmt_2100/return__
      -- CP-element group 78: 	 branch_block_stmt_2100/assign_stmt_2466__exit__
      -- CP-element group 78: 	 branch_block_stmt_2100/branch_block_stmt_2100__exit__
      -- CP-element group 78: 	 branch_block_stmt_2100/$exit
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2100/merge_stmt_2468_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2100/assign_stmt_2466/WPIPE_Block2_done_2463_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2100/assign_stmt_2466/$exit
      -- CP-element group 78: 	 branch_block_stmt_2100/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2100/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2100/merge_stmt_2468_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2100/merge_stmt_2468_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2100/merge_stmt_2468_PhiAck/dummy
      -- 
    ack_6185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2463_inst_ack_1, ack => convTransposeC_CP_5505_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_req
      -- CP-element group 79: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2237_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2233/$exit
      -- CP-element group 79: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/$exit
      -- 
    phi_stmt_2233_req_6196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2233_req_6196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(79), ack => phi_stmt_2233_req_0); -- 
    -- Element group convTransposeC_CP_5505_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5505_elements(43), ack => convTransposeC_CP_5505_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2240/$exit
      -- CP-element group 80: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2244_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- 
    phi_stmt_2240_req_6204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_6204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(80), ack => phi_stmt_2240_req_0); -- 
    -- Element group convTransposeC_CP_5505_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5505_elements(43), ack => convTransposeC_CP_5505_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Sample/$exit
      -- 
    ra_6221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_0, ack => convTransposeC_CP_5505_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Update/ca
      -- CP-element group 82: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/Update/$exit
      -- 
    ca_6226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_1, ack => convTransposeC_CP_5505_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_req
      -- CP-element group 83: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/SplitProtocol/$exit
      -- CP-element group 83: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2252/$exit
      -- CP-element group 83: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2247/$exit
      -- 
    phi_stmt_2247_req_6227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2247_req_6227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(83), ack => phi_stmt_2247_req_1); -- 
    convTransposeC_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(81) & convTransposeC_CP_5505_elements(82);
      gj_convTransposeC_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2226/$exit
      -- CP-element group 84: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2230_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_req
      -- CP-element group 84: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/$exit
      -- 
    phi_stmt_2226_req_6235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2226_req_6235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(84), ack => phi_stmt_2226_req_0); -- 
    -- Element group convTransposeC_CP_5505_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeC_CP_5505_elements(43), ack => convTransposeC_CP_5505_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2100/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(79) & convTransposeC_CP_5505_elements(80) & convTransposeC_CP_5505_elements(83) & convTransposeC_CP_5505_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Sample/$exit
      -- 
    ra_6255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2239_inst_ack_0, ack => convTransposeC_CP_5505_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Update/ca
      -- CP-element group 87: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/Update/$exit
      -- 
    ca_6260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2239_inst_ack_1, ack => convTransposeC_CP_5505_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/type_cast_2239/$exit
      -- CP-element group 88: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/$exit
      -- CP-element group 88: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2233/phi_stmt_2233_req
      -- 
    phi_stmt_2233_req_6261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2233_req_6261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(88), ack => phi_stmt_2233_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(86) & convTransposeC_CP_5505_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/$exit
      -- 
    ra_6278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2246_inst_ack_0, ack => convTransposeC_CP_5505_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/ca
      -- 
    ca_6283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2246_inst_ack_1, ack => convTransposeC_CP_5505_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/$exit
      -- CP-element group 91: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- CP-element group 91: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/$exit
      -- 
    phi_stmt_2240_req_6284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_6284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(91), ack => phi_stmt_2240_req_1); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(89) & convTransposeC_CP_5505_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Sample/$exit
      -- 
    ra_6301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2250_inst_ack_0, ack => convTransposeC_CP_5505_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Update/ca
      -- CP-element group 93: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/Update/$exit
      -- 
    ca_6306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2250_inst_ack_1, ack => convTransposeC_CP_5505_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_req
      -- CP-element group 94: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2250/$exit
      -- CP-element group 94: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/$exit
      -- 
    phi_stmt_2247_req_6307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2247_req_6307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(94), ack => phi_stmt_2247_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(92) & convTransposeC_CP_5505_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Sample/$exit
      -- 
    ra_6324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2232_inst_ack_0, ack => convTransposeC_CP_5505_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/Update/ca
      -- 
    ca_6329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2232_inst_ack_1, ack => convTransposeC_CP_5505_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2232/$exit
      -- CP-element group 97: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_req
      -- CP-element group 97: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2226/$exit
      -- 
    phi_stmt_2226_req_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2226_req_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(97), ack => phi_stmt_2226_req_1); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(95) & convTransposeC_CP_5505_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2100/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(88) & convTransposeC_CP_5505_elements(91) & convTransposeC_CP_5505_elements(94) & convTransposeC_CP_5505_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2100/merge_stmt_2225_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2100/merge_stmt_2225_PhiAck/$entry
      -- 
    convTransposeC_CP_5505_elements(99) <= OrReduce(convTransposeC_CP_5505_elements(85) & convTransposeC_CP_5505_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2100/merge_stmt_2225_PhiAck/phi_stmt_2226_ack
      -- 
    phi_stmt_2226_ack_6335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2226_ack_0, ack => convTransposeC_CP_5505_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2100/merge_stmt_2225_PhiAck/phi_stmt_2233_ack
      -- 
    phi_stmt_2233_ack_6336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2233_ack_0, ack => convTransposeC_CP_5505_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2100/merge_stmt_2225_PhiAck/phi_stmt_2240_ack
      -- 
    phi_stmt_2240_ack_6337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2240_ack_0, ack => convTransposeC_CP_5505_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2100/merge_stmt_2225_PhiAck/phi_stmt_2247_ack
      -- 
    phi_stmt_2247_ack_6338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2247_ack_0, ack => convTransposeC_CP_5505_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375__entry__
      -- CP-element group 104: 	 branch_block_stmt_2100/merge_stmt_2225__exit__
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2354_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/merge_stmt_2225_PhiAck/$exit
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2358_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2363_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2287_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2291_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2295_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/type_cast_2325_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/array_obj_ref_2331_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2332_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/ptr_deref_2336_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2100/assign_stmt_2259_to_assign_stmt_2375/addr_of_2355_update_start_
      -- 
    cr_6078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => ptr_deref_2358_store_0_req_1); -- 
    req_6013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => array_obj_ref_2354_index_offset_req_1); -- 
    cr_6092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2363_inst_req_1); -- 
    rr_6087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2363_inst_req_0); -- 
    req_6028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => addr_of_2355_final_reg_req_1); -- 
    rr_5839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2287_inst_req_0); -- 
    cr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2287_inst_req_1); -- 
    rr_5853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2291_inst_req_0); -- 
    cr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2291_inst_req_1); -- 
    rr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2295_inst_req_0); -- 
    cr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2295_inst_req_1); -- 
    rr_5881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2325_inst_req_0); -- 
    cr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => type_cast_2325_inst_req_1); -- 
    req_5917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => array_obj_ref_2331_index_offset_req_1); -- 
    req_5932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => addr_of_2332_final_reg_req_1); -- 
    cr_5977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(104), ack => ptr_deref_2336_load_0_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(100) & convTransposeC_CP_5505_elements(101) & convTransposeC_CP_5505_elements(102) & convTransposeC_CP_5505_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2434/$exit
      -- CP-element group 105: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2440_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_req
      -- 
    phi_stmt_2434_req_6373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2434_req_6373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(105), ack => phi_stmt_2434_req_1); -- 
    -- Element group convTransposeC_CP_5505_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5505_elements(76), ack => convTransposeC_CP_5505_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Sample/ra
      -- 
    ra_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2444_inst_ack_0, ack => convTransposeC_CP_5505_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/Update/ca
      -- 
    ca_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2444_inst_ack_1, ack => convTransposeC_CP_5505_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/$exit
      -- CP-element group 108: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/$exit
      -- CP-element group 108: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2444/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_req
      -- 
    phi_stmt_2441_req_6396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2441_req_6396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(108), ack => phi_stmt_2441_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(106) & convTransposeC_CP_5505_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Sample/ra
      -- 
    ra_6413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_0, ack => convTransposeC_CP_5505_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/Update/ca
      -- 
    ca_6418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_1, ack => convTransposeC_CP_5505_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/$exit
      -- CP-element group 111: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/$exit
      -- CP-element group 111: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2450/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_req
      -- 
    phi_stmt_2447_req_6419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2447_req_6419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(111), ack => phi_stmt_2447_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(109) & convTransposeC_CP_5505_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2100/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(105) & convTransposeC_CP_5505_elements(108) & convTransposeC_CP_5505_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/ra
      -- 
    ra_6439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_0, ack => convTransposeC_CP_5505_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/ca
      -- 
    ca_6444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_1, ack => convTransposeC_CP_5505_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/$exit
      -- CP-element group 115: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/$exit
      -- CP-element group 115: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2434/phi_stmt_2434_req
      -- 
    phi_stmt_2434_req_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2434_req_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(115), ack => phi_stmt_2434_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(113) & convTransposeC_CP_5505_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Sample/ra
      -- 
    ra_6462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2446_inst_ack_0, ack => convTransposeC_CP_5505_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/Update/ca
      -- 
    ca_6467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2446_inst_ack_1, ack => convTransposeC_CP_5505_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/$exit
      -- CP-element group 118: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/$exit
      -- CP-element group 118: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_sources/type_cast_2446/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2441/phi_stmt_2441_req
      -- 
    phi_stmt_2441_req_6468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2441_req_6468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(118), ack => phi_stmt_2441_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(116) & convTransposeC_CP_5505_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Sample/ra
      -- 
    ra_6485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2452_inst_ack_0, ack => convTransposeC_CP_5505_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/Update/ca
      -- 
    ca_6490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2452_inst_ack_1, ack => convTransposeC_CP_5505_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/$exit
      -- CP-element group 121: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/$exit
      -- CP-element group 121: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_sources/type_cast_2452/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2447/phi_stmt_2447_req
      -- 
    phi_stmt_2447_req_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2447_req_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5505_elements(121), ack => phi_stmt_2447_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(119) & convTransposeC_CP_5505_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2100/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(115) & convTransposeC_CP_5505_elements(118) & convTransposeC_CP_5505_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2100/merge_stmt_2433_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2100/merge_stmt_2433_PhiAck/$entry
      -- 
    convTransposeC_CP_5505_elements(123) <= OrReduce(convTransposeC_CP_5505_elements(112) & convTransposeC_CP_5505_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2100/merge_stmt_2433_PhiAck/phi_stmt_2434_ack
      -- 
    phi_stmt_2434_ack_6496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2434_ack_0, ack => convTransposeC_CP_5505_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2100/merge_stmt_2433_PhiAck/phi_stmt_2441_ack
      -- 
    phi_stmt_2441_ack_6497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2441_ack_0, ack => convTransposeC_CP_5505_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2100/merge_stmt_2433_PhiAck/phi_stmt_2447_ack
      -- 
    phi_stmt_2447_ack_6498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2447_ack_0, ack => convTransposeC_CP_5505_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2100/merge_stmt_2433_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5505_elements(124) & convTransposeC_CP_5505_elements(125) & convTransposeC_CP_5505_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5505_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2353_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2353_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2330_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2330_scaled : std_logic_vector(13 downto 0);
    signal add121_2223 : std_logic_vector(31 downto 0);
    signal add45_2174 : std_logic_vector(15 downto 0);
    signal add58_2185 : std_logic_vector(15 downto 0);
    signal add77_2306 : std_logic_vector(63 downto 0);
    signal add79_2316 : std_logic_vector(63 downto 0);
    signal add91_2370 : std_logic_vector(31 downto 0);
    signal add98_2388 : std_logic_vector(15 downto 0);
    signal add_2152 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2264 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2331_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2331_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2331_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2331_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2331_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2331_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2354_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2354_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2354_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2354_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2354_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2354_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2333 : std_logic_vector(31 downto 0);
    signal arrayidx87_2356 : std_logic_vector(31 downto 0);
    signal call11_2121 : std_logic_vector(15 downto 0);
    signal call13_2124 : std_logic_vector(15 downto 0);
    signal call14_2127 : std_logic_vector(15 downto 0);
    signal call15_2130 : std_logic_vector(15 downto 0);
    signal call16_2143 : std_logic_vector(15 downto 0);
    signal call18_2155 : std_logic_vector(15 downto 0);
    signal call1_2106 : std_logic_vector(15 downto 0);
    signal call20_2158 : std_logic_vector(15 downto 0);
    signal call22_2161 : std_logic_vector(15 downto 0);
    signal call3_2109 : std_logic_vector(15 downto 0);
    signal call5_2112 : std_logic_vector(15 downto 0);
    signal call7_2115 : std_logic_vector(15 downto 0);
    signal call9_2118 : std_logic_vector(15 downto 0);
    signal call_2103 : std_logic_vector(15 downto 0);
    signal cmp106_2401 : std_logic_vector(0 downto 0);
    signal cmp122_2426 : std_logic_vector(0 downto 0);
    signal cmp_2375 : std_logic_vector(0 downto 0);
    signal conv112_2421 : std_logic_vector(31 downto 0);
    signal conv115_2206 : std_logic_vector(31 downto 0);
    signal conv17_2147 : std_logic_vector(31 downto 0);
    signal conv65_2288 : std_logic_vector(63 downto 0);
    signal conv68_2194 : std_logic_vector(63 downto 0);
    signal conv70_2292 : std_logic_vector(63 downto 0);
    signal conv73_2198 : std_logic_vector(63 downto 0);
    signal conv75_2296 : std_logic_vector(63 downto 0);
    signal conv90_2364 : std_logic_vector(31 downto 0);
    signal conv94_2202 : std_logic_vector(31 downto 0);
    signal conv_2134 : std_logic_vector(31 downto 0);
    signal idxprom86_2349 : std_logic_vector(63 downto 0);
    signal idxprom_2326 : std_logic_vector(63 downto 0);
    signal inc110_2405 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2410 : std_logic_vector(15 downto 0);
    signal inc_2396 : std_logic_vector(15 downto 0);
    signal indvar_2226 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2459 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2447 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2247 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2441 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2240 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2417 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2434 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2233 : std_logic_vector(15 downto 0);
    signal mul54_2279 : std_logic_vector(15 downto 0);
    signal mul76_2301 : std_logic_vector(63 downto 0);
    signal mul78_2311 : std_logic_vector(63 downto 0);
    signal mul_2269 : std_logic_vector(15 downto 0);
    signal ptr_deref_2336_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2336_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2336_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2336_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2336_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2358_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2358_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2358_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2358_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2358_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2358_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2140 : std_logic_vector(31 downto 0);
    signal shr116137_2212 : std_logic_vector(31 downto 0);
    signal shr120138_2218 : std_logic_vector(31 downto 0);
    signal shr136_2168 : std_logic_vector(15 downto 0);
    signal shr81_2322 : std_logic_vector(31 downto 0);
    signal shr85_2343 : std_logic_vector(63 downto 0);
    signal sub48_2274 : std_logic_vector(15 downto 0);
    signal sub61_2190 : std_logic_vector(15 downto 0);
    signal sub62_2284 : std_logic_vector(15 downto 0);
    signal sub_2179 : std_logic_vector(15 downto 0);
    signal tmp1_2259 : std_logic_vector(31 downto 0);
    signal tmp83_2337 : std_logic_vector(63 downto 0);
    signal type_cast_2138_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2166_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2172_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2183_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2210_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2216_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2230_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2232_wire : std_logic_vector(31 downto 0);
    signal type_cast_2237_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2239_wire : std_logic_vector(15 downto 0);
    signal type_cast_2244_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2246_wire : std_logic_vector(15 downto 0);
    signal type_cast_2250_wire : std_logic_vector(15 downto 0);
    signal type_cast_2252_wire : std_logic_vector(15 downto 0);
    signal type_cast_2257_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2320_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2341_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2347_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2368_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2386_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2394_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2414_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2437_wire : std_logic_vector(15 downto 0);
    signal type_cast_2440_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2444_wire : std_logic_vector(15 downto 0);
    signal type_cast_2446_wire : std_logic_vector(15 downto 0);
    signal type_cast_2450_wire : std_logic_vector(15 downto 0);
    signal type_cast_2452_wire : std_logic_vector(15 downto 0);
    signal type_cast_2457_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2465_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2331_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2331_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2331_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2331_resized_base_address <= "00000000000000";
    array_obj_ref_2354_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2354_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2354_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2354_resized_base_address <= "00000000000000";
    ptr_deref_2336_word_offset_0 <= "00000000000000";
    ptr_deref_2358_word_offset_0 <= "00000000000000";
    type_cast_2138_wire_constant <= "00000000000000000000000000010000";
    type_cast_2166_wire_constant <= "0000000000000001";
    type_cast_2172_wire_constant <= "1111111111111111";
    type_cast_2183_wire_constant <= "1111111111111111";
    type_cast_2210_wire_constant <= "00000000000000000000000000000010";
    type_cast_2216_wire_constant <= "00000000000000000000000000000001";
    type_cast_2230_wire_constant <= "00000000000000000000000000000000";
    type_cast_2237_wire_constant <= "0000000000000000";
    type_cast_2244_wire_constant <= "0000000000000000";
    type_cast_2257_wire_constant <= "00000000000000000000000000000100";
    type_cast_2320_wire_constant <= "00000000000000000000000000000010";
    type_cast_2341_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2347_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2368_wire_constant <= "00000000000000000000000000000100";
    type_cast_2386_wire_constant <= "0000000000000100";
    type_cast_2394_wire_constant <= "0000000000000001";
    type_cast_2414_wire_constant <= "0000000000000000";
    type_cast_2440_wire_constant <= "0000000000000000";
    type_cast_2457_wire_constant <= "00000000000000000000000000000001";
    type_cast_2465_wire_constant <= "0000000000000001";
    phi_stmt_2226: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2230_wire_constant & type_cast_2232_wire;
      req <= phi_stmt_2226_req_0 & phi_stmt_2226_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2226",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2226_ack_0,
          idata => idata,
          odata => indvar_2226,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2226
    phi_stmt_2233: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2237_wire_constant & type_cast_2239_wire;
      req <= phi_stmt_2233_req_0 & phi_stmt_2233_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2233",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2233_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2233,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2233
    phi_stmt_2240: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2244_wire_constant & type_cast_2246_wire;
      req <= phi_stmt_2240_req_0 & phi_stmt_2240_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2240",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2240_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2240,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2240
    phi_stmt_2247: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2250_wire & type_cast_2252_wire;
      req <= phi_stmt_2247_req_0 & phi_stmt_2247_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2247",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2247_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2247,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2247
    phi_stmt_2434: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2437_wire & type_cast_2440_wire_constant;
      req <= phi_stmt_2434_req_0 & phi_stmt_2434_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2434",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2434_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2434,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2434
    phi_stmt_2441: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2444_wire & type_cast_2446_wire;
      req <= phi_stmt_2441_req_0 & phi_stmt_2441_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2441",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2441_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2441,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2441
    phi_stmt_2447: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2450_wire & type_cast_2452_wire;
      req <= phi_stmt_2447_req_0 & phi_stmt_2447_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2447",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2447_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2447,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2447
    -- flow-through select operator MUX_2416_inst
    input_dim1x_x2_2417 <= type_cast_2414_wire_constant when (cmp106_2401(0) /=  '0') else inc_2396;
    addr_of_2332_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2332_final_reg_req_0;
      addr_of_2332_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2332_final_reg_req_1;
      addr_of_2332_final_reg_ack_1<= rack(0);
      addr_of_2332_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2332_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2331_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2355_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2355_final_reg_req_0;
      addr_of_2355_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2355_final_reg_req_1;
      addr_of_2355_final_reg_ack_1<= rack(0);
      addr_of_2355_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2355_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2354_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2356,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2133_inst_req_0;
      type_cast_2133_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2133_inst_req_1;
      type_cast_2133_inst_ack_1<= rack(0);
      type_cast_2133_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2133_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2134,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2146_inst_req_0;
      type_cast_2146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2146_inst_req_1;
      type_cast_2146_inst_ack_1<= rack(0);
      type_cast_2146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2193_inst_req_0;
      type_cast_2193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2193_inst_req_1;
      type_cast_2193_inst_ack_1<= rack(0);
      type_cast_2193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2197_inst_req_0;
      type_cast_2197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2197_inst_req_1;
      type_cast_2197_inst_ack_1<= rack(0);
      type_cast_2197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2198,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2201_inst_req_0;
      type_cast_2201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2201_inst_req_1;
      type_cast_2201_inst_ack_1<= rack(0);
      type_cast_2201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2205_inst_req_0;
      type_cast_2205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2205_inst_req_1;
      type_cast_2205_inst_ack_1<= rack(0);
      type_cast_2205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2232_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2232_inst_req_0;
      type_cast_2232_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2232_inst_req_1;
      type_cast_2232_inst_ack_1<= rack(0);
      type_cast_2232_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2232_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2232_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2239_inst_req_0;
      type_cast_2239_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2239_inst_req_1;
      type_cast_2239_inst_ack_1<= rack(0);
      type_cast_2239_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2239_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2239_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2246_inst_req_0;
      type_cast_2246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2246_inst_req_1;
      type_cast_2246_inst_ack_1<= rack(0);
      type_cast_2246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2246_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2246_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2250_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2250_inst_req_0;
      type_cast_2250_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2250_inst_req_1;
      type_cast_2250_inst_ack_1<= rack(0);
      type_cast_2250_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2250_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2447,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2250_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2252_inst_req_0;
      type_cast_2252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2252_inst_req_1;
      type_cast_2252_inst_ack_1<= rack(0);
      type_cast_2252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2252_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2287_inst_req_0;
      type_cast_2287_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2287_inst_req_1;
      type_cast_2287_inst_ack_1<= rack(0);
      type_cast_2287_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2287_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2233,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2291_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2291_inst_req_0;
      type_cast_2291_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2291_inst_req_1;
      type_cast_2291_inst_ack_1<= rack(0);
      type_cast_2291_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2291_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2295_inst_req_0;
      type_cast_2295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2295_inst_req_1;
      type_cast_2295_inst_ack_1<= rack(0);
      type_cast_2295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2274,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2325_inst_req_0;
      type_cast_2325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2325_inst_req_1;
      type_cast_2325_inst_ack_1<= rack(0);
      type_cast_2325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2326,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2363_inst_req_0;
      type_cast_2363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2363_inst_req_1;
      type_cast_2363_inst_ack_1<= rack(0);
      type_cast_2363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2233,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2404_inst_req_0;
      type_cast_2404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2404_inst_req_1;
      type_cast_2404_inst_ack_1<= rack(0);
      type_cast_2404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2401,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2405,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2420_inst_req_0;
      type_cast_2420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2420_inst_req_1;
      type_cast_2420_inst_ack_1<= rack(0);
      type_cast_2420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2410,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2437_inst_req_0;
      type_cast_2437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2437_inst_req_1;
      type_cast_2437_inst_ack_1<= rack(0);
      type_cast_2437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2437_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2444_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2444_inst_req_0;
      type_cast_2444_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2444_inst_req_1;
      type_cast_2444_inst_ack_1<= rack(0);
      type_cast_2444_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2444_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2417,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2444_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2446_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2446_inst_req_0;
      type_cast_2446_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2446_inst_req_1;
      type_cast_2446_inst_ack_1<= rack(0);
      type_cast_2446_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2446_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2446_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2450_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2450_inst_req_0;
      type_cast_2450_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2450_inst_req_1;
      type_cast_2450_inst_ack_1<= rack(0);
      type_cast_2450_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2450_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2410,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2450_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2452_inst_req_0;
      type_cast_2452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2452_inst_req_1;
      type_cast_2452_inst_ack_1<= rack(0);
      type_cast_2452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2452_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2331_index_1_rename
    process(R_idxprom_2330_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2330_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2330_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2331_index_1_resize
    process(idxprom_2326) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2326;
      ov := iv(13 downto 0);
      R_idxprom_2330_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2331_root_address_inst
    process(array_obj_ref_2331_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2331_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2331_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2354_index_1_rename
    process(R_idxprom86_2353_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2353_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2353_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2354_index_1_resize
    process(idxprom86_2349) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2349;
      ov := iv(13 downto 0);
      R_idxprom86_2353_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2354_root_address_inst
    process(array_obj_ref_2354_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2354_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2354_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2336_addr_0
    process(ptr_deref_2336_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2336_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2336_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2336_base_resize
    process(arrayidx82_2333) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2333;
      ov := iv(13 downto 0);
      ptr_deref_2336_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2336_gather_scatter
    process(ptr_deref_2336_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2336_data_0;
      ov(63 downto 0) := iv;
      tmp83_2337 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2336_root_address_inst
    process(ptr_deref_2336_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2336_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2336_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_addr_0
    process(ptr_deref_2358_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2358_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_base_resize
    process(arrayidx87_2356) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2356;
      ov := iv(13 downto 0);
      ptr_deref_2358_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_gather_scatter
    process(tmp83_2337) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2337;
      ov(63 downto 0) := iv;
      ptr_deref_2358_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_root_address_inst
    process(ptr_deref_2358_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2358_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2376_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2375;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2376_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2376_branch_req_0,
          ack0 => if_stmt_2376_branch_ack_0,
          ack1 => if_stmt_2376_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2427_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2426;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2427_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2427_branch_req_0,
          ack0 => if_stmt_2427_branch_ack_0,
          ack1 => if_stmt_2427_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2173_inst
    process(call7_2115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2115, type_cast_2172_wire_constant, tmp_var);
      add45_2174 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2184_inst
    process(call9_2118) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2118, type_cast_2183_wire_constant, tmp_var);
      add58_2185 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2273_inst
    process(sub_2179, mul_2269) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2179, mul_2269, tmp_var);
      sub48_2274 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2283_inst
    process(sub61_2190, mul54_2279) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2190, mul54_2279, tmp_var);
      sub62_2284 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2387_inst
    process(input_dim2x_x1_2233) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2233, type_cast_2386_wire_constant, tmp_var);
      add98_2388 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2395_inst
    process(input_dim1x_x1_2240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2240, type_cast_2394_wire_constant, tmp_var);
      inc_2396 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2409_inst
    process(inc110_2405, input_dim0x_x2_2247) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2405, input_dim0x_x2_2247, tmp_var);
      inc110x_xinput_dim0x_x2_2410 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2222_inst
    process(shr116137_2212, shr120138_2218) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2212, shr120138_2218, tmp_var);
      add121_2223 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2263_inst
    process(add_2152, tmp1_2259) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2152, tmp1_2259, tmp_var);
      add_src_0x_x0_2264 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2369_inst
    process(conv90_2364) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2364, type_cast_2368_wire_constant, tmp_var);
      add91_2370 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2458_inst
    process(indvar_2226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2226, type_cast_2457_wire_constant, tmp_var);
      indvarx_xnext_2459 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2305_inst
    process(mul76_2301, conv70_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2301, conv70_2292, tmp_var);
      add77_2306 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2315_inst
    process(mul78_2311, conv65_2288) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2311, conv65_2288, tmp_var);
      add79_2316 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2348_inst
    process(shr85_2343) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2343, type_cast_2347_wire_constant, tmp_var);
      idxprom86_2349 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2400_inst
    process(inc_2396, call1_2106) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2396, call1_2106, tmp_var);
      cmp106_2401 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2425_inst
    process(conv112_2421, add121_2223) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2421, add121_2223, tmp_var);
      cmp122_2426 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2167_inst
    process(call_2103) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2103, type_cast_2166_wire_constant, tmp_var);
      shr136_2168 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2211_inst
    process(conv115_2206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2206, type_cast_2210_wire_constant, tmp_var);
      shr116137_2212 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2217_inst
    process(conv115_2206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2206, type_cast_2216_wire_constant, tmp_var);
      shr120138_2218 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2321_inst
    process(add_src_0x_x0_2264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2264, type_cast_2320_wire_constant, tmp_var);
      shr81_2322 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2342_inst
    process(add79_2316) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2316, type_cast_2341_wire_constant, tmp_var);
      shr85_2343 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2268_inst
    process(input_dim0x_x2_2247, call13_2124) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2247, call13_2124, tmp_var);
      mul_2269 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2278_inst
    process(input_dim1x_x1_2240, call13_2124) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2240, call13_2124, tmp_var);
      mul54_2279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2258_inst
    process(indvar_2226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2226, type_cast_2257_wire_constant, tmp_var);
      tmp1_2259 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2300_inst
    process(conv75_2296, conv73_2198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2296, conv73_2198, tmp_var);
      mul76_2301 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2310_inst
    process(add77_2306, conv68_2194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2306, conv68_2194, tmp_var);
      mul78_2311 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2151_inst
    process(shl_2140, conv17_2147) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2140, conv17_2147, tmp_var);
      add_2152 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2139_inst
    process(conv_2134) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2134, type_cast_2138_wire_constant, tmp_var);
      shl_2140 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2178_inst
    process(add45_2174, call14_2127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2174, call14_2127, tmp_var);
      sub_2179 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2189_inst
    process(add58_2185, call14_2127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2185, call14_2127, tmp_var);
      sub61_2190 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2374_inst
    process(add91_2370, conv94_2202) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2370, conv94_2202, tmp_var);
      cmp_2375 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2331_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2330_scaled;
      array_obj_ref_2331_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2331_index_offset_req_0;
      array_obj_ref_2331_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2331_index_offset_req_1;
      array_obj_ref_2331_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2354_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2353_scaled;
      array_obj_ref_2354_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2354_index_offset_req_0;
      array_obj_ref_2354_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2354_index_offset_req_1;
      array_obj_ref_2354_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2336_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2336_load_0_req_0;
      ptr_deref_2336_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2336_load_0_req_1;
      ptr_deref_2336_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2336_word_address_0;
      ptr_deref_2336_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2358_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2358_store_0_req_0;
      ptr_deref_2358_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2358_store_0_req_1;
      ptr_deref_2358_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2358_word_address_0;
      data_in <= ptr_deref_2358_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2102_inst RPIPE_Block2_start_2105_inst RPIPE_Block2_start_2108_inst RPIPE_Block2_start_2111_inst RPIPE_Block2_start_2114_inst RPIPE_Block2_start_2117_inst RPIPE_Block2_start_2120_inst RPIPE_Block2_start_2123_inst RPIPE_Block2_start_2126_inst RPIPE_Block2_start_2129_inst RPIPE_Block2_start_2142_inst RPIPE_Block2_start_2154_inst RPIPE_Block2_start_2157_inst RPIPE_Block2_start_2160_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2102_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2105_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2108_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2111_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2114_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2117_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2120_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2123_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2126_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2129_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2142_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2154_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2157_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2160_inst_req_0;
      RPIPE_Block2_start_2102_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2105_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2108_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2111_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2114_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2117_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2120_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2123_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2126_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2129_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2142_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2154_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2157_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2160_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2102_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2105_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2108_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2111_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2114_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2117_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2120_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2123_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2126_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2129_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2142_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2154_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2157_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2160_inst_req_1;
      RPIPE_Block2_start_2102_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2105_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2108_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2111_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2114_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2117_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2120_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2123_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2126_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2129_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2142_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2154_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2157_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2160_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2103 <= data_out(223 downto 208);
      call1_2106 <= data_out(207 downto 192);
      call3_2109 <= data_out(191 downto 176);
      call5_2112 <= data_out(175 downto 160);
      call7_2115 <= data_out(159 downto 144);
      call9_2118 <= data_out(143 downto 128);
      call11_2121 <= data_out(127 downto 112);
      call13_2124 <= data_out(111 downto 96);
      call14_2127 <= data_out(95 downto 80);
      call15_2130 <= data_out(79 downto 64);
      call16_2143 <= data_out(63 downto 48);
      call18_2155 <= data_out(47 downto 32);
      call20_2158 <= data_out(31 downto 16);
      call22_2161 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2463_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2463_inst_req_0;
      WPIPE_Block2_done_2463_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2463_inst_req_1;
      WPIPE_Block2_done_2463_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2465_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6515_start: Boolean;
  signal convTransposeD_CP_6515_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2483_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2483_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2480_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2477_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2483_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2480_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2480_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2477_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2477_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2480_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2483_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2486_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2486_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2486_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2486_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2492_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2492_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2498_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2492_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2498_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2495_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2498_inst_ack_1 : boolean;
  signal type_cast_2804_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2495_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2495_inst_ack_0 : boolean;
  signal if_stmt_2785_branch_ack_0 : boolean;
  signal RPIPE_Block3_start_2495_inst_req_0 : boolean;
  signal type_cast_2804_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2492_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2498_inst_req_0 : boolean;
  signal type_cast_2612_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2489_inst_req_0 : boolean;
  signal type_cast_2505_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2501_inst_req_1 : boolean;
  signal type_cast_2608_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2501_inst_ack_1 : boolean;
  signal phi_stmt_2799_req_0 : boolean;
  signal RPIPE_Block3_start_2501_inst_req_0 : boolean;
  signal type_cast_2608_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2501_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2477_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2474_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2474_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2489_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2489_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2474_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2474_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2489_inst_ack_0 : boolean;
  signal type_cast_2612_inst_ack_0 : boolean;
  signal type_cast_2808_inst_req_1 : boolean;
  signal type_cast_2808_inst_ack_1 : boolean;
  signal phi_stmt_2799_req_1 : boolean;
  signal type_cast_2802_inst_req_0 : boolean;
  signal type_cast_2591_inst_req_0 : boolean;
  signal type_cast_2591_inst_ack_0 : boolean;
  signal type_cast_2612_inst_req_1 : boolean;
  signal type_cast_2612_inst_ack_1 : boolean;
  signal type_cast_2802_inst_ack_0 : boolean;
  signal type_cast_2802_inst_req_1 : boolean;
  signal phi_stmt_2609_req_0 : boolean;
  signal type_cast_2808_inst_ack_0 : boolean;
  signal type_cast_2802_inst_ack_1 : boolean;
  signal phi_stmt_2805_req_0 : boolean;
  signal if_stmt_2785_branch_req_0 : boolean;
  signal type_cast_2608_inst_req_1 : boolean;
  signal type_cast_2591_inst_req_1 : boolean;
  signal type_cast_2505_inst_ack_0 : boolean;
  signal type_cast_2505_inst_req_1 : boolean;
  signal type_cast_2505_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2514_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2514_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2514_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2514_inst_ack_1 : boolean;
  signal type_cast_2518_inst_req_0 : boolean;
  signal type_cast_2518_inst_ack_0 : boolean;
  signal type_cast_2518_inst_req_1 : boolean;
  signal type_cast_2518_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2526_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2526_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2526_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2526_inst_ack_1 : boolean;
  signal if_stmt_2738_branch_ack_0 : boolean;
  signal RPIPE_Block3_start_2529_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2529_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2529_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2529_inst_ack_1 : boolean;
  signal phi_stmt_2805_req_1 : boolean;
  signal RPIPE_Block3_start_2532_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2532_inst_ack_0 : boolean;
  signal type_cast_2766_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2532_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2532_inst_ack_1 : boolean;
  signal type_cast_2810_inst_ack_1 : boolean;
  signal type_cast_2810_inst_req_1 : boolean;
  signal type_cast_2810_inst_ack_0 : boolean;
  signal phi_stmt_2602_req_0 : boolean;
  signal type_cast_2810_inst_req_0 : boolean;
  signal phi_stmt_2609_ack_0 : boolean;
  signal type_cast_2576_inst_req_0 : boolean;
  signal type_cast_2576_inst_ack_0 : boolean;
  signal type_cast_2804_inst_ack_0 : boolean;
  signal type_cast_2804_inst_req_0 : boolean;
  signal type_cast_2576_inst_req_1 : boolean;
  signal type_cast_2576_inst_ack_1 : boolean;
  signal phi_stmt_2792_req_0 : boolean;
  signal phi_stmt_2602_ack_0 : boolean;
  signal phi_stmt_2595_ack_0 : boolean;
  signal type_cast_2580_inst_req_0 : boolean;
  signal type_cast_2580_inst_ack_0 : boolean;
  signal type_cast_2580_inst_req_1 : boolean;
  signal type_cast_2580_inst_ack_1 : boolean;
  signal type_cast_2795_inst_ack_1 : boolean;
  signal type_cast_2795_inst_req_1 : boolean;
  signal phi_stmt_2588_ack_0 : boolean;
  signal type_cast_2584_inst_req_0 : boolean;
  signal type_cast_2584_inst_ack_0 : boolean;
  signal type_cast_2584_inst_req_1 : boolean;
  signal phi_stmt_2595_req_1 : boolean;
  signal type_cast_2584_inst_ack_1 : boolean;
  signal phi_stmt_2609_req_1 : boolean;
  signal type_cast_2601_inst_ack_1 : boolean;
  signal type_cast_2649_inst_req_0 : boolean;
  signal type_cast_2649_inst_ack_0 : boolean;
  signal type_cast_2601_inst_req_1 : boolean;
  signal type_cast_2649_inst_req_1 : boolean;
  signal type_cast_2649_inst_ack_1 : boolean;
  signal if_stmt_2738_branch_ack_1 : boolean;
  signal type_cast_2795_inst_ack_0 : boolean;
  signal type_cast_2614_inst_ack_1 : boolean;
  signal type_cast_2614_inst_req_1 : boolean;
  signal type_cast_2653_inst_req_0 : boolean;
  signal type_cast_2653_inst_ack_0 : boolean;
  signal type_cast_2653_inst_req_1 : boolean;
  signal type_cast_2653_inst_ack_1 : boolean;
  signal type_cast_2795_inst_req_0 : boolean;
  signal type_cast_2614_inst_ack_0 : boolean;
  signal type_cast_2657_inst_req_0 : boolean;
  signal type_cast_2601_inst_ack_0 : boolean;
  signal type_cast_2657_inst_ack_0 : boolean;
  signal type_cast_2657_inst_req_1 : boolean;
  signal type_cast_2601_inst_req_0 : boolean;
  signal type_cast_2657_inst_ack_1 : boolean;
  signal type_cast_2614_inst_req_0 : boolean;
  signal phi_stmt_2595_req_0 : boolean;
  signal type_cast_2687_inst_req_0 : boolean;
  signal type_cast_2687_inst_ack_0 : boolean;
  signal type_cast_2687_inst_req_1 : boolean;
  signal type_cast_2687_inst_ack_1 : boolean;
  signal type_cast_2808_inst_req_0 : boolean;
  signal phi_stmt_2792_req_1 : boolean;
  signal phi_stmt_2588_req_1 : boolean;
  signal array_obj_ref_2693_index_offset_req_0 : boolean;
  signal array_obj_ref_2693_index_offset_ack_0 : boolean;
  signal type_cast_2766_inst_req_1 : boolean;
  signal array_obj_ref_2693_index_offset_req_1 : boolean;
  signal array_obj_ref_2693_index_offset_ack_1 : boolean;
  signal addr_of_2694_final_reg_req_0 : boolean;
  signal addr_of_2694_final_reg_ack_0 : boolean;
  signal if_stmt_2738_branch_req_0 : boolean;
  signal addr_of_2694_final_reg_req_1 : boolean;
  signal addr_of_2694_final_reg_ack_1 : boolean;
  signal type_cast_2766_inst_ack_0 : boolean;
  signal phi_stmt_2602_req_1 : boolean;
  signal WPIPE_Block3_done_2821_inst_ack_1 : boolean;
  signal type_cast_2766_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2821_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2821_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2821_inst_req_0 : boolean;
  signal phi_stmt_2588_req_0 : boolean;
  signal if_stmt_2785_branch_ack_1 : boolean;
  signal ptr_deref_2698_load_0_req_0 : boolean;
  signal ptr_deref_2698_load_0_ack_0 : boolean;
  signal ptr_deref_2698_load_0_req_1 : boolean;
  signal ptr_deref_2698_load_0_ack_1 : boolean;
  signal type_cast_2591_inst_ack_1 : boolean;
  signal type_cast_2608_inst_ack_1 : boolean;
  signal array_obj_ref_2716_index_offset_req_0 : boolean;
  signal array_obj_ref_2716_index_offset_ack_0 : boolean;
  signal array_obj_ref_2716_index_offset_req_1 : boolean;
  signal array_obj_ref_2716_index_offset_ack_1 : boolean;
  signal addr_of_2717_final_reg_req_0 : boolean;
  signal addr_of_2717_final_reg_ack_0 : boolean;
  signal addr_of_2717_final_reg_req_1 : boolean;
  signal addr_of_2717_final_reg_ack_1 : boolean;
  signal ptr_deref_2720_store_0_req_0 : boolean;
  signal ptr_deref_2720_store_0_ack_0 : boolean;
  signal ptr_deref_2720_store_0_req_1 : boolean;
  signal ptr_deref_2720_store_0_ack_1 : boolean;
  signal type_cast_2725_inst_req_0 : boolean;
  signal type_cast_2725_inst_ack_0 : boolean;
  signal type_cast_2725_inst_req_1 : boolean;
  signal type_cast_2725_inst_ack_1 : boolean;
  signal phi_stmt_2792_ack_0 : boolean;
  signal phi_stmt_2799_ack_0 : boolean;
  signal phi_stmt_2805_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6515_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6515_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6515_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6515_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6515: Block -- control-path 
    signal convTransposeD_CP_6515_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6515_elements(0) <= convTransposeD_CP_6515_start;
    convTransposeD_CP_6515_symbol <= convTransposeD_CP_6515_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2472/$entry
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/$entry
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533__entry__
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2472/branch_block_stmt_2472__entry__
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Update/cr
      -- 
    rr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(0), ack => RPIPE_Block3_start_2474_inst_req_0); -- 
    cr_6708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(0), ack => type_cast_2505_inst_req_1); -- 
    cr_6736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(0), ack => type_cast_2518_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2472/assign_stmt_2817/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2472/assign_stmt_2817__exit__
      -- CP-element group 1: 	 branch_block_stmt_2472/assign_stmt_2817__entry__
      -- CP-element group 1: 	 branch_block_stmt_2472/merge_stmt_2791__exit__
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/assign_stmt_2817/$exit
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/$entry
      -- CP-element group 1: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/$entry
      -- 
    rr_7282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2608_inst_req_0); -- 
    rr_7236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2591_inst_req_0); -- 
    cr_7287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2608_inst_req_1); -- 
    cr_7241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2591_inst_req_1); -- 
    cr_7264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2601_inst_req_1); -- 
    cr_7310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2614_inst_req_1); -- 
    rr_7259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2601_inst_req_0); -- 
    rr_7305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(1), ack => type_cast_2614_inst_req_0); -- 
    convTransposeD_CP_6515_elements(1) <= convTransposeD_CP_6515_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Sample/$exit
      -- 
    ra_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2474_inst_ack_0, ack => convTransposeD_CP_6515_elements(2)); -- 
    cr_6568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(2), ack => RPIPE_Block3_start_2474_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2474_Update/$exit
      -- 
    ca_6569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2474_inst_ack_1, ack => convTransposeD_CP_6515_elements(3)); -- 
    rr_6577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(3), ack => RPIPE_Block3_start_2477_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_sample_completed_
      -- 
    ra_6578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2477_inst_ack_0, ack => convTransposeD_CP_6515_elements(4)); -- 
    cr_6582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(4), ack => RPIPE_Block3_start_2477_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2477_update_completed_
      -- 
    ca_6583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2477_inst_ack_1, ack => convTransposeD_CP_6515_elements(5)); -- 
    rr_6591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(5), ack => RPIPE_Block3_start_2480_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_sample_completed_
      -- 
    ra_6592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2480_inst_ack_0, ack => convTransposeD_CP_6515_elements(6)); -- 
    cr_6596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(6), ack => RPIPE_Block3_start_2480_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2480_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Sample/$entry
      -- 
    ca_6597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2480_inst_ack_1, ack => convTransposeD_CP_6515_elements(7)); -- 
    rr_6605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(7), ack => RPIPE_Block3_start_2483_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Sample/$exit
      -- 
    ra_6606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2483_inst_ack_0, ack => convTransposeD_CP_6515_elements(8)); -- 
    cr_6610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(8), ack => RPIPE_Block3_start_2483_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2483_update_completed_
      -- 
    ca_6611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2483_inst_ack_1, ack => convTransposeD_CP_6515_elements(9)); -- 
    rr_6619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(9), ack => RPIPE_Block3_start_2486_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_sample_completed_
      -- 
    ra_6620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2486_inst_ack_0, ack => convTransposeD_CP_6515_elements(10)); -- 
    cr_6624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(10), ack => RPIPE_Block3_start_2486_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2486_update_completed_
      -- 
    ca_6625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2486_inst_ack_1, ack => convTransposeD_CP_6515_elements(11)); -- 
    rr_6633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(11), ack => RPIPE_Block3_start_2489_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Sample/ra
      -- 
    ra_6634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2489_inst_ack_0, ack => convTransposeD_CP_6515_elements(12)); -- 
    cr_6638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(12), ack => RPIPE_Block3_start_2489_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2489_Update/$exit
      -- 
    ca_6639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2489_inst_ack_1, ack => convTransposeD_CP_6515_elements(13)); -- 
    rr_6647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(13), ack => RPIPE_Block3_start_2492_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_sample_completed_
      -- 
    ra_6648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2492_inst_ack_0, ack => convTransposeD_CP_6515_elements(14)); -- 
    cr_6652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(14), ack => RPIPE_Block3_start_2492_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2492_update_completed_
      -- 
    ca_6653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2492_inst_ack_1, ack => convTransposeD_CP_6515_elements(15)); -- 
    rr_6661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(15), ack => RPIPE_Block3_start_2495_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_sample_completed_
      -- 
    ra_6662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2495_inst_ack_0, ack => convTransposeD_CP_6515_elements(16)); -- 
    cr_6666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(16), ack => RPIPE_Block3_start_2495_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2495_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Sample/rr
      -- 
    ca_6667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2495_inst_ack_1, ack => convTransposeD_CP_6515_elements(17)); -- 
    rr_6675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(17), ack => RPIPE_Block3_start_2498_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Sample/ra
      -- 
    ra_6676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2498_inst_ack_0, ack => convTransposeD_CP_6515_elements(18)); -- 
    cr_6680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(18), ack => RPIPE_Block3_start_2498_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2498_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Sample/$entry
      -- 
    ca_6681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2498_inst_ack_1, ack => convTransposeD_CP_6515_elements(19)); -- 
    rr_6689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(19), ack => RPIPE_Block3_start_2501_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_update_start_
      -- 
    ra_6690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2501_inst_ack_0, ack => convTransposeD_CP_6515_elements(20)); -- 
    cr_6694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(20), ack => RPIPE_Block3_start_2501_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2501_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Sample/rr
      -- 
    ca_6695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2501_inst_ack_1, ack => convTransposeD_CP_6515_elements(21)); -- 
    rr_6703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(21), ack => type_cast_2505_inst_req_0); -- 
    rr_6717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(21), ack => RPIPE_Block3_start_2514_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Sample/ra
      -- 
    ra_6704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2505_inst_ack_0, ack => convTransposeD_CP_6515_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2505_Update/ca
      -- 
    ca_6709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2505_inst_ack_1, ack => convTransposeD_CP_6515_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Update/cr
      -- 
    ra_6718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2514_inst_ack_0, ack => convTransposeD_CP_6515_elements(24)); -- 
    cr_6722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(24), ack => RPIPE_Block3_start_2514_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2514_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Sample/rr
      -- 
    ca_6723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2514_inst_ack_1, ack => convTransposeD_CP_6515_elements(25)); -- 
    rr_6731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(25), ack => type_cast_2518_inst_req_0); -- 
    rr_6745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(25), ack => RPIPE_Block3_start_2526_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Sample/ra
      -- 
    ra_6732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_0, ack => convTransposeD_CP_6515_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/type_cast_2518_Update/ca
      -- 
    ca_6737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_1, ack => convTransposeD_CP_6515_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Update/cr
      -- 
    ra_6746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2526_inst_ack_0, ack => convTransposeD_CP_6515_elements(28)); -- 
    cr_6750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(28), ack => RPIPE_Block3_start_2526_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2526_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Sample/rr
      -- 
    ca_6751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2526_inst_ack_1, ack => convTransposeD_CP_6515_elements(29)); -- 
    rr_6759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(29), ack => RPIPE_Block3_start_2529_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Update/cr
      -- 
    ra_6760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2529_inst_ack_0, ack => convTransposeD_CP_6515_elements(30)); -- 
    cr_6764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(30), ack => RPIPE_Block3_start_2529_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2529_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Sample/rr
      -- 
    ca_6765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2529_inst_ack_1, ack => convTransposeD_CP_6515_elements(31)); -- 
    rr_6773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(31), ack => RPIPE_Block3_start_2532_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Update/cr
      -- 
    ra_6774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2532_inst_ack_0, ack => convTransposeD_CP_6515_elements(32)); -- 
    cr_6778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(32), ack => RPIPE_Block3_start_2532_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/RPIPE_Block3_start_2532_Update/ca
      -- 
    ca_6779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2532_inst_ack_1, ack => convTransposeD_CP_6515_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533/$exit
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585__entry__
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2475_to_assign_stmt_2533__exit__
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/$entry
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Update/cr
      -- 
    rr_6790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(34), ack => type_cast_2576_inst_req_0); -- 
    cr_6795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(34), ack => type_cast_2576_inst_req_1); -- 
    rr_6804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(34), ack => type_cast_2580_inst_req_0); -- 
    cr_6809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(34), ack => type_cast_2580_inst_req_1); -- 
    rr_6818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(34), ack => type_cast_2584_inst_req_0); -- 
    cr_6823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(34), ack => type_cast_2584_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(23) & convTransposeD_CP_6515_elements(27) & convTransposeD_CP_6515_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Sample/ra
      -- 
    ra_6791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2576_inst_ack_0, ack => convTransposeD_CP_6515_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2576_Update/ca
      -- 
    ca_6796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2576_inst_ack_1, ack => convTransposeD_CP_6515_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Sample/ra
      -- 
    ra_6805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2580_inst_ack_0, ack => convTransposeD_CP_6515_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2580_Update/ca
      -- 
    ca_6810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2580_inst_ack_1, ack => convTransposeD_CP_6515_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Sample/ra
      -- 
    ra_6819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2584_inst_ack_0, ack => convTransposeD_CP_6515_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/type_cast_2584_Update/ca
      -- 
    ca_6824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2584_inst_ack_1, ack => convTransposeD_CP_6515_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585__exit__
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/assign_stmt_2540_to_assign_stmt_2585/$exit
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2602/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2595/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2588/$entry
      -- CP-element group 41: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/$entry
      -- 
    rr_7210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(41), ack => type_cast_2612_inst_req_0); -- 
    cr_7215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(41), ack => type_cast_2612_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(36) & convTransposeD_CP_6515_elements(38) & convTransposeD_CP_6515_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Sample/ra
      -- 
    ra_6836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2649_inst_ack_0, ack => convTransposeD_CP_6515_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Update/ca
      -- 
    ca_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2649_inst_ack_1, ack => convTransposeD_CP_6515_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Sample/ra
      -- 
    ra_6850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2653_inst_ack_0, ack => convTransposeD_CP_6515_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Update/ca
      -- 
    ca_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2653_inst_ack_1, ack => convTransposeD_CP_6515_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Sample/ra
      -- 
    ra_6864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2657_inst_ack_0, ack => convTransposeD_CP_6515_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Update/ca
      -- 
    ca_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2657_inst_ack_1, ack => convTransposeD_CP_6515_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Sample/ra
      -- 
    ra_6878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2687_inst_ack_0, ack => convTransposeD_CP_6515_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Sample/req
      -- 
    ca_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2687_inst_ack_1, ack => convTransposeD_CP_6515_elements(49)); -- 
    req_6908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(49), ack => array_obj_ref_2693_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Sample/ack
      -- 
    ack_6909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2693_index_offset_ack_0, ack => convTransposeD_CP_6515_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_request/req
      -- 
    ack_6914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2693_index_offset_ack_1, ack => convTransposeD_CP_6515_elements(51)); -- 
    req_6923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(51), ack => addr_of_2694_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_request/ack
      -- 
    ack_6924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2694_final_reg_ack_0, ack => convTransposeD_CP_6515_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/word_access_start/word_0/rr
      -- 
    ack_6929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2694_final_reg_ack_1, ack => convTransposeD_CP_6515_elements(53)); -- 
    rr_6962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(53), ack => ptr_deref_2698_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Sample/word_access_start/word_0/ra
      -- 
    ra_6963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2698_load_0_ack_0, ack => convTransposeD_CP_6515_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/ptr_deref_2698_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/ptr_deref_2698_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/ptr_deref_2698_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/ptr_deref_2698_Merge/merge_ack
      -- 
    ca_6974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2698_load_0_ack_1, ack => convTransposeD_CP_6515_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Sample/req
      -- 
    req_7004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(56), ack => array_obj_ref_2716_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(43) & convTransposeD_CP_6515_elements(45) & convTransposeD_CP_6515_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Sample/ack
      -- 
    ack_7005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2716_index_offset_ack_0, ack => convTransposeD_CP_6515_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_request/req
      -- 
    ack_7010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2716_index_offset_ack_1, ack => convTransposeD_CP_6515_elements(58)); -- 
    req_7019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(58), ack => addr_of_2717_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_request/ack
      -- 
    ack_7020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2717_final_reg_ack_0, ack => convTransposeD_CP_6515_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_word_addrgen/root_register_ack
      -- 
    ack_7025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2717_final_reg_ack_1, ack => convTransposeD_CP_6515_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/ptr_deref_2720_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/ptr_deref_2720_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/ptr_deref_2720_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/ptr_deref_2720_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/word_access_start/word_0/rr
      -- 
    rr_7063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(61), ack => ptr_deref_2720_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(55) & convTransposeD_CP_6515_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Sample/word_access_start/word_0/ra
      -- 
    ra_7064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2720_store_0_ack_0, ack => convTransposeD_CP_6515_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/word_access_complete/word_0/ca
      -- 
    ca_7075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2720_store_0_ack_1, ack => convTransposeD_CP_6515_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Sample/ra
      -- 
    ra_7084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2725_inst_ack_0, ack => convTransposeD_CP_6515_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Update/ca
      -- 
    ca_7089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2725_inst_ack_1, ack => convTransposeD_CP_6515_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737__exit__
      -- CP-element group 66: 	 branch_block_stmt_2472/if_stmt_2738__entry__
      -- CP-element group 66: 	 branch_block_stmt_2472/if_stmt_2738_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/$exit
      -- CP-element group 66: 	 branch_block_stmt_2472/if_stmt_2738_else_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2472/R_cmp_2739_place
      -- CP-element group 66: 	 branch_block_stmt_2472/if_stmt_2738_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2472/if_stmt_2738_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2472/if_stmt_2738_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2472/if_stmt_2738_dead_link/$entry
      -- 
    branch_req_7097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(66), ack => if_stmt_2738_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(50) & convTransposeD_CP_6515_elements(57) & convTransposeD_CP_6515_elements(63) & convTransposeD_CP_6515_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2472/merge_stmt_2744__exit__
      -- CP-element group 67: 	 branch_block_stmt_2472/assign_stmt_2750__entry__
      -- CP-element group 67: 	 branch_block_stmt_2472/assign_stmt_2750__exit__
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2472/merge_stmt_2744_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2472/merge_stmt_2744_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2472/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/merge_stmt_2744_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2472/merge_stmt_2744_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2472/if_stmt_2738_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/assign_stmt_2750/$exit
      -- CP-element group 67: 	 branch_block_stmt_2472/assign_stmt_2750/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/if_stmt_2738_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2472/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Sample/rr
      -- 
    if_choice_transition_7102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2738_branch_ack_1, ack => convTransposeD_CP_6515_elements(67)); -- 
    cr_7471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(67), ack => type_cast_2808_inst_req_1); -- 
    rr_7443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(67), ack => type_cast_2802_inst_req_0); -- 
    cr_7448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(67), ack => type_cast_2802_inst_req_1); -- 
    cr_7425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(67), ack => type_cast_2795_inst_req_1); -- 
    rr_7420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(67), ack => type_cast_2795_inst_req_0); -- 
    rr_7466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(67), ack => type_cast_2808_inst_req_0); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784__entry__
      -- CP-element group 68: 	 branch_block_stmt_2472/merge_stmt_2752__exit__
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2472/merge_stmt_2752_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2472/merge_stmt_2752_PhiAck/dummy
      -- CP-element group 68: 	 branch_block_stmt_2472/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2472/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2472/merge_stmt_2752_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2472/merge_stmt_2752_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/$entry
      -- CP-element group 68: 	 branch_block_stmt_2472/if_stmt_2738_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2472/if_stmt_2738_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2472/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Sample/$entry
      -- 
    else_choice_transition_7106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2738_branch_ack_0, ack => convTransposeD_CP_6515_elements(68)); -- 
    cr_7127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(68), ack => type_cast_2766_inst_req_1); -- 
    rr_7122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(68), ack => type_cast_2766_inst_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Sample/$exit
      -- 
    ra_7123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_0, ack => convTransposeD_CP_6515_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2472/if_stmt_2785__entry__
      -- CP-element group 70: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784__exit__
      -- CP-element group 70: 	 branch_block_stmt_2472/if_stmt_2785_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2472/if_stmt_2785_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2472/if_stmt_2785_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/$exit
      -- CP-element group 70: 	 branch_block_stmt_2472/if_stmt_2785_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2472/R_cmp121_2786_place
      -- CP-element group 70: 	 branch_block_stmt_2472/if_stmt_2785_else_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2472/assign_stmt_2758_to_assign_stmt_2784/type_cast_2766_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2472/if_stmt_2785_if_link/$entry
      -- 
    ca_7128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_1, ack => convTransposeD_CP_6515_elements(70)); -- 
    branch_req_7136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(70), ack => if_stmt_2785_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2472/assign_stmt_2824__entry__
      -- CP-element group 71: 	 branch_block_stmt_2472/merge_stmt_2819__exit__
      -- CP-element group 71: 	 branch_block_stmt_2472/assign_stmt_2824/$entry
      -- CP-element group 71: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2472/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2472/if_stmt_2785_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2472/if_stmt_2785_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2472/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2472/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2472/merge_stmt_2819_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2472/merge_stmt_2819_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2472/merge_stmt_2819_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2472/merge_stmt_2819_PhiAck/dummy
      -- 
    if_choice_transition_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2785_branch_ack_1, ack => convTransposeD_CP_6515_elements(71)); -- 
    req_7161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(71), ack => WPIPE_Block3_done_2821_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2472/if_stmt_2785_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2472/if_stmt_2785_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2792/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/$entry
      -- CP-element group 72: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/$entry
      -- 
    else_choice_transition_7145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2785_branch_ack_0, ack => convTransposeD_CP_6515_elements(72)); -- 
    cr_7376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(72), ack => type_cast_2804_inst_req_1); -- 
    cr_7399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(72), ack => type_cast_2810_inst_req_1); -- 
    rr_7394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(72), ack => type_cast_2810_inst_req_0); -- 
    rr_7371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(72), ack => type_cast_2804_inst_req_0); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Update/req
      -- CP-element group 73: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Sample/$exit
      -- 
    ack_7162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2821_inst_ack_0, ack => convTransposeD_CP_6515_elements(73)); -- 
    req_7166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(73), ack => WPIPE_Block3_done_2821_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2472/$exit
      -- CP-element group 74: 	 branch_block_stmt_2472/merge_stmt_2826__exit__
      -- CP-element group 74: 	 branch_block_stmt_2472/return__
      -- CP-element group 74: 	 branch_block_stmt_2472/assign_stmt_2824__exit__
      -- CP-element group 74: 	 branch_block_stmt_2472/branch_block_stmt_2472__exit__
      -- CP-element group 74: 	 branch_block_stmt_2472/assign_stmt_2824/$exit
      -- CP-element group 74: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2472/assign_stmt_2824/WPIPE_Block3_done_2821_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2472/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2472/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2472/merge_stmt_2826_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2472/merge_stmt_2826_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2472/merge_stmt_2826_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2472/merge_stmt_2826_PhiAck/dummy
      -- 
    ack_7167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2821_inst_ack_1, ack => convTransposeD_CP_6515_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_req
      -- CP-element group 75: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2594_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2588/$exit
      -- 
    phi_stmt_2588_req_7178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2588_req_7178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(75), ack => phi_stmt_2588_req_1); -- 
    -- Element group convTransposeD_CP_6515_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6515_elements(41), ack => convTransposeD_CP_6515_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_req
      -- CP-element group 76: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2599_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2595/$exit
      -- 
    phi_stmt_2595_req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2595_req_7186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(76), ack => phi_stmt_2595_req_0); -- 
    -- Element group convTransposeD_CP_6515_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6515_elements(41), ack => convTransposeD_CP_6515_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_req
      -- CP-element group 77: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2606_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2602/$exit
      -- 
    phi_stmt_2602_req_7194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2602_req_7194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(77), ack => phi_stmt_2602_req_0); -- 
    -- Element group convTransposeD_CP_6515_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6515_elements(41), ack => convTransposeD_CP_6515_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Sample/ra
      -- 
    ra_7211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2612_inst_ack_0, ack => convTransposeD_CP_6515_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/Update/ca
      -- 
    ca_7216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2612_inst_ack_1, ack => convTransposeD_CP_6515_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2612/$exit
      -- CP-element group 80: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_req
      -- CP-element group 80: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/phi_stmt_2609/$exit
      -- 
    phi_stmt_2609_req_7217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2609_req_7217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(80), ack => phi_stmt_2609_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(78) & convTransposeD_CP_6515_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2472/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(75) & convTransposeD_CP_6515_elements(76) & convTransposeD_CP_6515_elements(77) & convTransposeD_CP_6515_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Sample/ra
      -- 
    ra_7237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2591_inst_ack_0, ack => convTransposeD_CP_6515_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/Update/ca
      -- 
    ca_7242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2591_inst_ack_1, ack => convTransposeD_CP_6515_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/$exit
      -- CP-element group 84: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_sources/type_cast_2591/$exit
      -- CP-element group 84: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2588/phi_stmt_2588_req
      -- 
    phi_stmt_2588_req_7243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2588_req_7243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(84), ack => phi_stmt_2588_req_0); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(82) & convTransposeD_CP_6515_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Sample/$exit
      -- 
    ra_7260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2601_inst_ack_0, ack => convTransposeD_CP_6515_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/Update/$exit
      -- 
    ca_7265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2601_inst_ack_1, ack => convTransposeD_CP_6515_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_req
      -- CP-element group 87: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2601/$exit
      -- CP-element group 87: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2595/$exit
      -- 
    phi_stmt_2595_req_7266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2595_req_7266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(87), ack => phi_stmt_2595_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(85) & convTransposeD_CP_6515_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/$exit
      -- 
    ra_7283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2608_inst_ack_0, ack => convTransposeD_CP_6515_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/ca
      -- 
    ca_7288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2608_inst_ack_1, ack => convTransposeD_CP_6515_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/$exit
      -- CP-element group 90: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/$exit
      -- CP-element group 90: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_req
      -- 
    phi_stmt_2602_req_7289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2602_req_7289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(90), ack => phi_stmt_2602_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(88) & convTransposeD_CP_6515_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Sample/$exit
      -- 
    ra_7306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_0, ack => convTransposeD_CP_6515_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Update/ca
      -- CP-element group 92: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/Update/$exit
      -- 
    ca_7311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_1, ack => convTransposeD_CP_6515_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_req
      -- CP-element group 93: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2614/$exit
      -- CP-element group 93: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/$exit
      -- 
    phi_stmt_2609_req_7312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2609_req_7312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(93), ack => phi_stmt_2609_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(91) & convTransposeD_CP_6515_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2472/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(84) & convTransposeD_CP_6515_elements(87) & convTransposeD_CP_6515_elements(90) & convTransposeD_CP_6515_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2472/merge_stmt_2587_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2472/merge_stmt_2587_PhiAck/$entry
      -- 
    convTransposeD_CP_6515_elements(95) <= OrReduce(convTransposeD_CP_6515_elements(81) & convTransposeD_CP_6515_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2472/merge_stmt_2587_PhiAck/phi_stmt_2588_ack
      -- 
    phi_stmt_2588_ack_7317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2588_ack_0, ack => convTransposeD_CP_6515_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2472/merge_stmt_2587_PhiAck/phi_stmt_2595_ack
      -- 
    phi_stmt_2595_ack_7318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2595_ack_0, ack => convTransposeD_CP_6515_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2472/merge_stmt_2587_PhiAck/phi_stmt_2602_ack
      -- 
    phi_stmt_2602_ack_7319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2602_ack_0, ack => convTransposeD_CP_6515_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2472/merge_stmt_2587_PhiAck/phi_stmt_2609_ack
      -- 
    phi_stmt_2609_ack_7320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2609_ack_0, ack => convTransposeD_CP_6515_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737__entry__
      -- CP-element group 100: 	 branch_block_stmt_2472/merge_stmt_2587__exit__
      -- CP-element group 100: 	 branch_block_stmt_2472/merge_stmt_2587_PhiAck/$exit
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2649_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2653_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2657_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2687_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2693_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2694_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2698_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/array_obj_ref_2716_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/addr_of_2717_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/ptr_deref_2720_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2472/assign_stmt_2621_to_assign_stmt_2737/type_cast_2725_Update/cr
      -- 
    rr_6835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2649_inst_req_0); -- 
    cr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2649_inst_req_1); -- 
    rr_6849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2653_inst_req_0); -- 
    cr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2653_inst_req_1); -- 
    rr_6863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2657_inst_req_0); -- 
    cr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2657_inst_req_1); -- 
    rr_6877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2687_inst_req_0); -- 
    cr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2687_inst_req_1); -- 
    req_6913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => array_obj_ref_2693_index_offset_req_1); -- 
    req_6928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => addr_of_2694_final_reg_req_1); -- 
    cr_6973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => ptr_deref_2698_load_0_req_1); -- 
    req_7009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => array_obj_ref_2716_index_offset_req_1); -- 
    req_7024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => addr_of_2717_final_reg_req_1); -- 
    cr_7074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => ptr_deref_2720_store_0_req_1); -- 
    rr_7083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2725_inst_req_0); -- 
    cr_7088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(100), ack => type_cast_2725_inst_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(96) & convTransposeD_CP_6515_elements(97) & convTransposeD_CP_6515_elements(98) & convTransposeD_CP_6515_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2792/$exit
      -- CP-element group 101: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_req
      -- CP-element group 101: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2798_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/$exit
      -- 
    phi_stmt_2792_req_7355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2792_req_7355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(101), ack => phi_stmt_2792_req_1); -- 
    -- Element group convTransposeD_CP_6515_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6515_elements(72), ack => convTransposeD_CP_6515_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/$exit
      -- 
    ra_7372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2804_inst_ack_0, ack => convTransposeD_CP_6515_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/ca
      -- CP-element group 103: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/$exit
      -- 
    ca_7377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2804_inst_ack_1, ack => convTransposeD_CP_6515_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_req
      -- CP-element group 104: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/$exit
      -- CP-element group 104: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2799/$exit
      -- 
    phi_stmt_2799_req_7378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2799_req_7378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(104), ack => phi_stmt_2799_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(102) & convTransposeD_CP_6515_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Sample/$exit
      -- 
    ra_7395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2810_inst_ack_0, ack => convTransposeD_CP_6515_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/Update/$exit
      -- 
    ca_7400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2810_inst_ack_1, ack => convTransposeD_CP_6515_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/$exit
      -- CP-element group 107: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_req
      -- CP-element group 107: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2810/$exit
      -- CP-element group 107: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/$exit
      -- 
    phi_stmt_2805_req_7401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2805_req_7401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(107), ack => phi_stmt_2805_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(105) & convTransposeD_CP_6515_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2472/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(101) & convTransposeD_CP_6515_elements(104) & convTransposeD_CP_6515_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Sample/$exit
      -- 
    ra_7421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2795_inst_ack_0, ack => convTransposeD_CP_6515_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Update/ca
      -- CP-element group 110: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/Update/$exit
      -- 
    ca_7426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2795_inst_ack_1, ack => convTransposeD_CP_6515_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/$exit
      -- CP-element group 111: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_req
      -- CP-element group 111: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2792/phi_stmt_2792_sources/type_cast_2795/$exit
      -- 
    phi_stmt_2792_req_7427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2792_req_7427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(111), ack => phi_stmt_2792_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(109) & convTransposeD_CP_6515_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/$exit
      -- 
    ra_7444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_0, ack => convTransposeD_CP_6515_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/ca
      -- 
    ca_7449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_1, ack => convTransposeD_CP_6515_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_req
      -- CP-element group 114: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/$exit
      -- CP-element group 114: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2799/$exit
      -- 
    phi_stmt_2799_req_7450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2799_req_7450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(114), ack => phi_stmt_2799_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(112) & convTransposeD_CP_6515_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Sample/ra
      -- 
    ra_7467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2808_inst_ack_0, ack => convTransposeD_CP_6515_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Update/ca
      -- CP-element group 116: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/Update/$exit
      -- 
    ca_7472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2808_inst_ack_1, ack => convTransposeD_CP_6515_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/$exit
      -- CP-element group 117: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_req
      -- CP-element group 117: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2805/phi_stmt_2805_sources/type_cast_2808/$exit
      -- 
    phi_stmt_2805_req_7473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2805_req_7473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6515_elements(117), ack => phi_stmt_2805_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(115) & convTransposeD_CP_6515_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2472/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(111) & convTransposeD_CP_6515_elements(114) & convTransposeD_CP_6515_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2472/merge_stmt_2791_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2472/merge_stmt_2791_PhiAck/$entry
      -- 
    convTransposeD_CP_6515_elements(119) <= OrReduce(convTransposeD_CP_6515_elements(108) & convTransposeD_CP_6515_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2472/merge_stmt_2791_PhiAck/phi_stmt_2792_ack
      -- 
    phi_stmt_2792_ack_7478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2792_ack_0, ack => convTransposeD_CP_6515_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2472/merge_stmt_2791_PhiAck/phi_stmt_2799_ack
      -- 
    phi_stmt_2799_ack_7479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2799_ack_0, ack => convTransposeD_CP_6515_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2472/merge_stmt_2791_PhiAck/phi_stmt_2805_ack
      -- 
    phi_stmt_2805_ack_7480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2805_ack_0, ack => convTransposeD_CP_6515_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2472/merge_stmt_2791_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6515_elements(120) & convTransposeD_CP_6515_elements(121) & convTransposeD_CP_6515_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6515_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2715_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2715_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2692_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2692_scaled : std_logic_vector(13 downto 0);
    signal add103_2750 : std_logic_vector(15 downto 0);
    signal add32_2551 : std_logic_vector(15 downto 0);
    signal add50_2557 : std_logic_vector(15 downto 0);
    signal add63_2568 : std_logic_vector(15 downto 0);
    signal add82_2668 : std_logic_vector(63 downto 0);
    signal add84_2678 : std_logic_vector(63 downto 0);
    signal add96_2732 : std_logic_vector(31 downto 0);
    signal add_2524 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2626 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2693_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2693_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2693_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2693_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2693_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2693_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2716_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2716_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2716_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2716_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2716_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2716_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2695 : std_logic_vector(31 downto 0);
    signal arrayidx92_2718 : std_logic_vector(31 downto 0);
    signal call11_2493 : std_logic_vector(15 downto 0);
    signal call13_2496 : std_logic_vector(15 downto 0);
    signal call14_2499 : std_logic_vector(15 downto 0);
    signal call15_2502 : std_logic_vector(15 downto 0);
    signal call16_2515 : std_logic_vector(15 downto 0);
    signal call18_2527 : std_logic_vector(15 downto 0);
    signal call1_2478 : std_logic_vector(15 downto 0);
    signal call20_2530 : std_logic_vector(15 downto 0);
    signal call22_2533 : std_logic_vector(15 downto 0);
    signal call3_2481 : std_logic_vector(15 downto 0);
    signal call5_2484 : std_logic_vector(15 downto 0);
    signal call7_2487 : std_logic_vector(15 downto 0);
    signal call9_2490 : std_logic_vector(15 downto 0);
    signal call_2475 : std_logic_vector(15 downto 0);
    signal cmp111_2763 : std_logic_vector(0 downto 0);
    signal cmp121_2784 : std_logic_vector(0 downto 0);
    signal cmp_2737 : std_logic_vector(0 downto 0);
    signal conv17_2519 : std_logic_vector(31 downto 0);
    signal conv70_2650 : std_logic_vector(63 downto 0);
    signal conv73_2577 : std_logic_vector(63 downto 0);
    signal conv75_2654 : std_logic_vector(63 downto 0);
    signal conv78_2581 : std_logic_vector(63 downto 0);
    signal conv80_2658 : std_logic_vector(63 downto 0);
    signal conv95_2726 : std_logic_vector(31 downto 0);
    signal conv99_2585 : std_logic_vector(31 downto 0);
    signal conv_2506 : std_logic_vector(31 downto 0);
    signal idxprom91_2711 : std_logic_vector(63 downto 0);
    signal idxprom_2688 : std_logic_vector(63 downto 0);
    signal inc115_2767 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2772 : std_logic_vector(15 downto 0);
    signal inc_2758 : std_logic_vector(15 downto 0);
    signal indvar_2588 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2817 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2805 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2609 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2799 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2602 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2779 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2792 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2595 : std_logic_vector(15 downto 0);
    signal mul59_2641 : std_logic_vector(15 downto 0);
    signal mul81_2663 : std_logic_vector(63 downto 0);
    signal mul83_2673 : std_logic_vector(63 downto 0);
    signal mul_2631 : std_logic_vector(15 downto 0);
    signal ptr_deref_2698_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2698_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2698_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2698_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2698_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2720_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2720_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2720_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2720_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2720_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2720_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2512 : std_logic_vector(31 downto 0);
    signal shr135_2540 : std_logic_vector(15 downto 0);
    signal shr31136_2546 : std_logic_vector(15 downto 0);
    signal shr86_2684 : std_logic_vector(31 downto 0);
    signal shr90_2705 : std_logic_vector(63 downto 0);
    signal sub53_2636 : std_logic_vector(15 downto 0);
    signal sub66_2573 : std_logic_vector(15 downto 0);
    signal sub67_2646 : std_logic_vector(15 downto 0);
    signal sub_2562 : std_logic_vector(15 downto 0);
    signal tmp1_2621 : std_logic_vector(31 downto 0);
    signal tmp88_2699 : std_logic_vector(63 downto 0);
    signal type_cast_2510_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2538_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2544_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2555_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2591_wire : std_logic_vector(31 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2599_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2601_wire : std_logic_vector(15 downto 0);
    signal type_cast_2606_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2608_wire : std_logic_vector(15 downto 0);
    signal type_cast_2612_wire : std_logic_vector(15 downto 0);
    signal type_cast_2614_wire : std_logic_vector(15 downto 0);
    signal type_cast_2619_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2682_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2703_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2709_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2730_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2748_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2756_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2776_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2795_wire : std_logic_vector(15 downto 0);
    signal type_cast_2798_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2802_wire : std_logic_vector(15 downto 0);
    signal type_cast_2804_wire : std_logic_vector(15 downto 0);
    signal type_cast_2808_wire : std_logic_vector(15 downto 0);
    signal type_cast_2810_wire : std_logic_vector(15 downto 0);
    signal type_cast_2815_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2823_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2693_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2693_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2693_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2693_resized_base_address <= "00000000000000";
    array_obj_ref_2716_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2716_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2716_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2716_resized_base_address <= "00000000000000";
    ptr_deref_2698_word_offset_0 <= "00000000000000";
    ptr_deref_2720_word_offset_0 <= "00000000000000";
    type_cast_2510_wire_constant <= "00000000000000000000000000010000";
    type_cast_2538_wire_constant <= "0000000000000010";
    type_cast_2544_wire_constant <= "0000000000000001";
    type_cast_2555_wire_constant <= "1111111111111111";
    type_cast_2566_wire_constant <= "1111111111111111";
    type_cast_2594_wire_constant <= "00000000000000000000000000000000";
    type_cast_2599_wire_constant <= "0000000000000000";
    type_cast_2606_wire_constant <= "0000000000000000";
    type_cast_2619_wire_constant <= "00000000000000000000000000000100";
    type_cast_2682_wire_constant <= "00000000000000000000000000000010";
    type_cast_2703_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2709_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2730_wire_constant <= "00000000000000000000000000000100";
    type_cast_2748_wire_constant <= "0000000000000100";
    type_cast_2756_wire_constant <= "0000000000000001";
    type_cast_2776_wire_constant <= "0000000000000000";
    type_cast_2798_wire_constant <= "0000000000000000";
    type_cast_2815_wire_constant <= "00000000000000000000000000000001";
    type_cast_2823_wire_constant <= "0000000000000001";
    phi_stmt_2588: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2591_wire & type_cast_2594_wire_constant;
      req <= phi_stmt_2588_req_0 & phi_stmt_2588_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2588",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2588_ack_0,
          idata => idata,
          odata => indvar_2588,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2588
    phi_stmt_2595: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2599_wire_constant & type_cast_2601_wire;
      req <= phi_stmt_2595_req_0 & phi_stmt_2595_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2595",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2595_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2595,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2595
    phi_stmt_2602: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2606_wire_constant & type_cast_2608_wire;
      req <= phi_stmt_2602_req_0 & phi_stmt_2602_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2602",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2602_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2602,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2602
    phi_stmt_2609: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2612_wire & type_cast_2614_wire;
      req <= phi_stmt_2609_req_0 & phi_stmt_2609_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2609",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2609_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2609,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2609
    phi_stmt_2792: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2795_wire & type_cast_2798_wire_constant;
      req <= phi_stmt_2792_req_0 & phi_stmt_2792_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2792",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2792_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2792,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2792
    phi_stmt_2799: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2802_wire & type_cast_2804_wire;
      req <= phi_stmt_2799_req_0 & phi_stmt_2799_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2799",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2799_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2799,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2799
    phi_stmt_2805: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2808_wire & type_cast_2810_wire;
      req <= phi_stmt_2805_req_0 & phi_stmt_2805_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2805",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2805_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2805,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2805
    -- flow-through select operator MUX_2778_inst
    input_dim1x_x2_2779 <= type_cast_2776_wire_constant when (cmp111_2763(0) /=  '0') else inc_2758;
    addr_of_2694_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2694_final_reg_req_0;
      addr_of_2694_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2694_final_reg_req_1;
      addr_of_2694_final_reg_ack_1<= rack(0);
      addr_of_2694_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2694_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2693_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2717_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2717_final_reg_req_0;
      addr_of_2717_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2717_final_reg_req_1;
      addr_of_2717_final_reg_ack_1<= rack(0);
      addr_of_2717_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2717_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2716_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2505_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2505_inst_req_0;
      type_cast_2505_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2505_inst_req_1;
      type_cast_2505_inst_ack_1<= rack(0);
      type_cast_2505_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2505_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2502,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2506,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2518_inst_req_0;
      type_cast_2518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2518_inst_req_1;
      type_cast_2518_inst_ack_1<= rack(0);
      type_cast_2518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2576_inst_req_0;
      type_cast_2576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2576_inst_req_1;
      type_cast_2576_inst_ack_1<= rack(0);
      type_cast_2576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2533,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2580_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2580_inst_req_0;
      type_cast_2580_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2580_inst_req_1;
      type_cast_2580_inst_ack_1<= rack(0);
      type_cast_2580_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2580_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2581,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2584_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2584_inst_req_0;
      type_cast_2584_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2584_inst_req_1;
      type_cast_2584_inst_ack_1<= rack(0);
      type_cast_2584_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2584_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2481,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2585,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2591_inst_req_0;
      type_cast_2591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2591_inst_req_1;
      type_cast_2591_inst_ack_1<= rack(0);
      type_cast_2591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2817,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2591_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2601_inst_req_0;
      type_cast_2601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2601_inst_req_1;
      type_cast_2601_inst_ack_1<= rack(0);
      type_cast_2601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2601_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2608_inst_req_0;
      type_cast_2608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2608_inst_req_1;
      type_cast_2608_inst_ack_1<= rack(0);
      type_cast_2608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2608_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2612_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2612_inst_req_0;
      type_cast_2612_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2612_inst_req_1;
      type_cast_2612_inst_ack_1<= rack(0);
      type_cast_2612_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2612_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2612_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2614_inst_req_0;
      type_cast_2614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2614_inst_req_1;
      type_cast_2614_inst_ack_1<= rack(0);
      type_cast_2614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2805,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2614_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2649_inst_req_0;
      type_cast_2649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2649_inst_req_1;
      type_cast_2649_inst_ack_1<= rack(0);
      type_cast_2649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2653_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2653_inst_req_0;
      type_cast_2653_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2653_inst_req_1;
      type_cast_2653_inst_ack_1<= rack(0);
      type_cast_2653_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2653_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2654,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2657_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2657_inst_req_0;
      type_cast_2657_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2657_inst_req_1;
      type_cast_2657_inst_ack_1<= rack(0);
      type_cast_2657_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2657_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2687_inst_req_0;
      type_cast_2687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2687_inst_req_1;
      type_cast_2687_inst_ack_1<= rack(0);
      type_cast_2687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2725_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2725_inst_req_0;
      type_cast_2725_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2725_inst_req_1;
      type_cast_2725_inst_ack_1<= rack(0);
      type_cast_2725_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2725_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2726,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2766_inst_req_0;
      type_cast_2766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2766_inst_req_1;
      type_cast_2766_inst_ack_1<= rack(0);
      type_cast_2766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2763,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2795_inst_req_0;
      type_cast_2795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2795_inst_req_1;
      type_cast_2795_inst_ack_1<= rack(0);
      type_cast_2795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2750,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2795_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2802_inst_req_0;
      type_cast_2802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2802_inst_req_1;
      type_cast_2802_inst_ack_1<= rack(0);
      type_cast_2802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2802_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2804_inst_req_0;
      type_cast_2804_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2804_inst_req_1;
      type_cast_2804_inst_ack_1<= rack(0);
      type_cast_2804_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2804_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2804_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2808_inst_req_0;
      type_cast_2808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2808_inst_req_1;
      type_cast_2808_inst_ack_1<= rack(0);
      type_cast_2808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2609,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2808_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2810_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2810_inst_req_0;
      type_cast_2810_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2810_inst_req_1;
      type_cast_2810_inst_ack_1<= rack(0);
      type_cast_2810_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2810_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2772,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2810_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2693_index_1_rename
    process(R_idxprom_2692_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2692_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2692_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2693_index_1_resize
    process(idxprom_2688) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2688;
      ov := iv(13 downto 0);
      R_idxprom_2692_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2693_root_address_inst
    process(array_obj_ref_2693_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2693_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2693_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2716_index_1_rename
    process(R_idxprom91_2715_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2715_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2715_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2716_index_1_resize
    process(idxprom91_2711) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2711;
      ov := iv(13 downto 0);
      R_idxprom91_2715_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2716_root_address_inst
    process(array_obj_ref_2716_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2716_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2716_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2698_addr_0
    process(ptr_deref_2698_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2698_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2698_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2698_base_resize
    process(arrayidx87_2695) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2695;
      ov := iv(13 downto 0);
      ptr_deref_2698_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2698_gather_scatter
    process(ptr_deref_2698_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2698_data_0;
      ov(63 downto 0) := iv;
      tmp88_2699 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2698_root_address_inst
    process(ptr_deref_2698_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2698_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2698_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2720_addr_0
    process(ptr_deref_2720_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2720_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2720_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2720_base_resize
    process(arrayidx92_2718) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2718;
      ov := iv(13 downto 0);
      ptr_deref_2720_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2720_gather_scatter
    process(tmp88_2699) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2699;
      ov(63 downto 0) := iv;
      ptr_deref_2720_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2720_root_address_inst
    process(ptr_deref_2720_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2720_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2720_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2738_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2737;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2738_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2738_branch_req_0,
          ack0 => if_stmt_2738_branch_ack_0,
          ack1 => if_stmt_2738_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2785_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2784;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2785_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2785_branch_req_0,
          ack0 => if_stmt_2785_branch_ack_0,
          ack1 => if_stmt_2785_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2550_inst
    process(shr135_2540, shr31136_2546) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2540, shr31136_2546, tmp_var);
      add32_2551 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2556_inst
    process(call7_2487) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2487, type_cast_2555_wire_constant, tmp_var);
      add50_2557 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2567_inst
    process(call9_2490) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2490, type_cast_2566_wire_constant, tmp_var);
      add63_2568 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2635_inst
    process(sub_2562, mul_2631) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2562, mul_2631, tmp_var);
      sub53_2636 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2645_inst
    process(sub66_2573, mul59_2641) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2573, mul59_2641, tmp_var);
      sub67_2646 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2749_inst
    process(input_dim2x_x1_2595) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2595, type_cast_2748_wire_constant, tmp_var);
      add103_2750 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2757_inst
    process(input_dim1x_x1_2602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2602, type_cast_2756_wire_constant, tmp_var);
      inc_2758 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2771_inst
    process(inc115_2767, input_dim0x_x2_2609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2767, input_dim0x_x2_2609, tmp_var);
      inc115x_xinput_dim0x_x2_2772 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2625_inst
    process(add_2524, tmp1_2621) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2524, tmp1_2621, tmp_var);
      add_src_0x_x0_2626 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2731_inst
    process(conv95_2726) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2726, type_cast_2730_wire_constant, tmp_var);
      add96_2732 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2816_inst
    process(indvar_2588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2588, type_cast_2815_wire_constant, tmp_var);
      indvarx_xnext_2817 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2667_inst
    process(mul81_2663, conv75_2654) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2663, conv75_2654, tmp_var);
      add82_2668 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2677_inst
    process(mul83_2673, conv70_2650) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2673, conv70_2650, tmp_var);
      add84_2678 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2710_inst
    process(shr90_2705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2705, type_cast_2709_wire_constant, tmp_var);
      idxprom91_2711 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2762_inst
    process(inc_2758, call1_2478) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2758, call1_2478, tmp_var);
      cmp111_2763 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2783_inst
    process(inc115x_xinput_dim0x_x2_2772, call_2475) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2772, call_2475, tmp_var);
      cmp121_2784 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2539_inst
    process(call_2475) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2475, type_cast_2538_wire_constant, tmp_var);
      shr135_2540 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2545_inst
    process(call_2475) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2475, type_cast_2544_wire_constant, tmp_var);
      shr31136_2546 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2683_inst
    process(add_src_0x_x0_2626) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2626, type_cast_2682_wire_constant, tmp_var);
      shr86_2684 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2704_inst
    process(add84_2678) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2678, type_cast_2703_wire_constant, tmp_var);
      shr90_2705 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2630_inst
    process(input_dim0x_x2_2609, call13_2496) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2609, call13_2496, tmp_var);
      mul_2631 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2640_inst
    process(input_dim1x_x1_2602, call13_2496) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2602, call13_2496, tmp_var);
      mul59_2641 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2620_inst
    process(indvar_2588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2588, type_cast_2619_wire_constant, tmp_var);
      tmp1_2621 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2662_inst
    process(conv80_2658, conv78_2581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2658, conv78_2581, tmp_var);
      mul81_2663 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2672_inst
    process(add82_2668, conv73_2577) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2668, conv73_2577, tmp_var);
      mul83_2673 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2523_inst
    process(shl_2512, conv17_2519) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2512, conv17_2519, tmp_var);
      add_2524 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2511_inst
    process(conv_2506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2506, type_cast_2510_wire_constant, tmp_var);
      shl_2512 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2561_inst
    process(add50_2557, call14_2499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2557, call14_2499, tmp_var);
      sub_2562 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2572_inst
    process(add63_2568, call14_2499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2568, call14_2499, tmp_var);
      sub66_2573 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2736_inst
    process(add96_2732, conv99_2585) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2732, conv99_2585, tmp_var);
      cmp_2737 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2693_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2692_scaled;
      array_obj_ref_2693_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2693_index_offset_req_0;
      array_obj_ref_2693_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2693_index_offset_req_1;
      array_obj_ref_2693_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2716_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2715_scaled;
      array_obj_ref_2716_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2716_index_offset_req_0;
      array_obj_ref_2716_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2716_index_offset_req_1;
      array_obj_ref_2716_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2698_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2698_load_0_req_0;
      ptr_deref_2698_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2698_load_0_req_1;
      ptr_deref_2698_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2698_word_address_0;
      ptr_deref_2698_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2720_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2720_store_0_req_0;
      ptr_deref_2720_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2720_store_0_req_1;
      ptr_deref_2720_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2720_word_address_0;
      data_in <= ptr_deref_2720_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2474_inst RPIPE_Block3_start_2477_inst RPIPE_Block3_start_2480_inst RPIPE_Block3_start_2483_inst RPIPE_Block3_start_2486_inst RPIPE_Block3_start_2489_inst RPIPE_Block3_start_2492_inst RPIPE_Block3_start_2495_inst RPIPE_Block3_start_2498_inst RPIPE_Block3_start_2501_inst RPIPE_Block3_start_2514_inst RPIPE_Block3_start_2526_inst RPIPE_Block3_start_2529_inst RPIPE_Block3_start_2532_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2474_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2477_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2480_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2483_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2486_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2489_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2492_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2495_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2498_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2501_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2514_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2526_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2529_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2532_inst_req_0;
      RPIPE_Block3_start_2474_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2477_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2480_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2483_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2486_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2489_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2492_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2495_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2498_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2501_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2514_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2526_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2529_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2532_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2474_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2477_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2480_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2483_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2486_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2489_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2492_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2495_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2498_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2501_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2514_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2526_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2529_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2532_inst_req_1;
      RPIPE_Block3_start_2474_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2477_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2480_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2483_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2486_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2489_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2492_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2495_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2498_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2501_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2514_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2526_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2529_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2532_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2475 <= data_out(223 downto 208);
      call1_2478 <= data_out(207 downto 192);
      call3_2481 <= data_out(191 downto 176);
      call5_2484 <= data_out(175 downto 160);
      call7_2487 <= data_out(159 downto 144);
      call9_2490 <= data_out(143 downto 128);
      call11_2493 <= data_out(127 downto 112);
      call13_2496 <= data_out(111 downto 96);
      call14_2499 <= data_out(95 downto 80);
      call15_2502 <= data_out(79 downto 64);
      call16_2515 <= data_out(63 downto 48);
      call18_2527 <= data_out(47 downto 32);
      call20_2530 <= data_out(31 downto 16);
      call22_2533 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2821_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2821_inst_req_0;
      WPIPE_Block3_done_2821_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2821_inst_req_1;
      WPIPE_Block3_done_2821_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2823_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(10 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(4 downto 4),
      memory_space_2_sr_ack => memory_space_2_sr_ack(4 downto 4),
      memory_space_2_sr_addr => memory_space_2_sr_addr(69 downto 56),
      memory_space_2_sr_data => memory_space_2_sr_data(319 downto 256),
      memory_space_2_sr_tag => memory_space_2_sr_tag(94 downto 76),
      memory_space_2_sc_req => memory_space_2_sc_req(4 downto 4),
      memory_space_2_sc_ack => memory_space_2_sc_ack(4 downto 4),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(55 downto 42),
      memory_space_0_lr_tag => memory_space_0_lr_tag(75 downto 57),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(255 downto 192),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 3),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 3),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 3),
      memory_space_2_sr_addr => memory_space_2_sr_addr(55 downto 42),
      memory_space_2_sr_data => memory_space_2_sr_data(255 downto 192),
      memory_space_2_sr_tag => memory_space_2_sr_tag(75 downto 57),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 3),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 3),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(41 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(56 downto 38),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(191 downto 128),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 2),
      memory_space_2_sr_req => memory_space_2_sr_req(2 downto 2),
      memory_space_2_sr_ack => memory_space_2_sr_ack(2 downto 2),
      memory_space_2_sr_addr => memory_space_2_sr_addr(41 downto 28),
      memory_space_2_sr_data => memory_space_2_sr_data(191 downto 128),
      memory_space_2_sr_tag => memory_space_2_sr_tag(56 downto 38),
      memory_space_2_sc_req => memory_space_2_sc_req(2 downto 2),
      memory_space_2_sc_ack => memory_space_2_sc_ack(2 downto 2),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 1),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(27 downto 14),
      memory_space_2_sr_data => memory_space_2_sr_data(127 downto 64),
      memory_space_2_sr_tag => memory_space_2_sr_tag(37 downto 19),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
