-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    ct_core_call_reqs : out  std_logic_vector(0 downto 0);
    ct_core_call_acks : in   std_logic_vector(0 downto 0);
    ct_core_call_data : out  std_logic_vector(175 downto 0);
    ct_core_call_tag  :  out  std_logic_vector(0 downto 0);
    ct_core_return_reqs : out  std_logic_vector(0 downto 0);
    ct_core_return_acks : in   std_logic_vector(0 downto 0);
    ct_core_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_772_start: Boolean;
  signal convTranspose_CP_772_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component ct_core is -- 
    generic (tag_length : integer); 
    port ( -- 
      inp_d0 : in  std_logic_vector(15 downto 0);
      inp_d1 : in  std_logic_vector(15 downto 0);
      inp_d2 : in  std_logic_vector(15 downto 0);
      ker_d1 : in  std_logic_vector(15 downto 0);
      ker_d2 : in  std_logic_vector(15 downto 0);
      out_d0 : in  std_logic_vector(15 downto 0);
      out_d1 : in  std_logic_vector(15 downto 0);
      out_d2 : in  std_logic_vector(15 downto 0);
      stride : in  std_logic_vector(15 downto 0);
      padding : in  std_logic_vector(15 downto 0);
      index1 : in  std_logic_vector(7 downto 0);
      index3 : in  std_logic_vector(7 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(39 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(0 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(103 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_data : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_ConvTranspose_input_pipe_477_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_464_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_377_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1528_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_427_inst_ack_1 : boolean;
  signal type_cast_1500_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_427_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_377_inst_req_1 : boolean;
  signal type_cast_800_inst_ack_1 : boolean;
  signal ptr_deref_880_store_0_req_1 : boolean;
  signal type_cast_481_inst_req_1 : boolean;
  signal type_cast_393_inst_ack_0 : boolean;
  signal type_cast_381_inst_ack_0 : boolean;
  signal type_cast_431_inst_req_0 : boolean;
  signal type_cast_393_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_850_inst_ack_0 : boolean;
  signal type_cast_431_inst_req_1 : boolean;
  signal type_cast_431_inst_ack_1 : boolean;
  signal type_cast_356_inst_req_1 : boolean;
  signal type_cast_998_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_389_inst_req_0 : boolean;
  signal type_cast_512_inst_req_0 : boolean;
  signal type_cast_481_inst_ack_0 : boolean;
  signal type_cast_498_inst_req_0 : boolean;
  signal type_cast_406_inst_req_0 : boolean;
  signal type_cast_980_inst_ack_1 : boolean;
  signal type_cast_468_inst_ack_0 : boolean;
  signal type_cast_443_inst_ack_0 : boolean;
  signal type_cast_800_inst_req_1 : boolean;
  signal type_cast_331_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_ack_0 : boolean;
  signal type_cast_980_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_452_inst_ack_1 : boolean;
  signal type_cast_381_inst_req_0 : boolean;
  signal type_cast_393_inst_req_0 : boolean;
  signal type_cast_1016_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_464_inst_req_1 : boolean;
  signal type_cast_381_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_339_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_req_0 : boolean;
  signal type_cast_331_inst_ack_1 : boolean;
  signal type_cast_406_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_452_inst_req_0 : boolean;
  signal type_cast_456_inst_req_1 : boolean;
  signal type_cast_418_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_339_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_439_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_389_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_377_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1364_inst_req_0 : boolean;
  signal type_cast_343_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_339_inst_req_0 : boolean;
  signal type_cast_418_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_439_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_ack_1 : boolean;
  signal type_cast_1034_inst_req_1 : boolean;
  signal type_cast_1016_inst_req_0 : boolean;
  signal type_cast_1016_inst_ack_0 : boolean;
  signal type_cast_490_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1030_inst_ack_1 : boolean;
  signal type_cast_512_inst_ack_0 : boolean;
  signal type_cast_494_inst_ack_1 : boolean;
  signal type_cast_356_inst_req_0 : boolean;
  signal type_cast_468_inst_req_0 : boolean;
  signal type_cast_356_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_452_inst_req_1 : boolean;
  signal type_cast_494_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_477_inst_ack_0 : boolean;
  signal type_cast_516_inst_req_1 : boolean;
  signal type_cast_516_inst_ack_1 : boolean;
  signal type_cast_443_inst_req_0 : boolean;
  signal array_obj_ref_959_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_389_inst_ack_0 : boolean;
  signal type_cast_443_inst_req_1 : boolean;
  signal addr_of_960_final_reg_req_0 : boolean;
  signal type_cast_494_inst_ack_0 : boolean;
  signal type_cast_998_inst_ack_0 : boolean;
  signal type_cast_331_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1084_inst_ack_1 : boolean;
  signal type_cast_481_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_389_inst_ack_1 : boolean;
  signal type_cast_406_inst_req_1 : boolean;
  signal type_cast_406_inst_ack_1 : boolean;
  signal type_cast_356_inst_ack_1 : boolean;
  signal type_cast_443_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_377_inst_ack_1 : boolean;
  signal type_cast_456_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_339_inst_ack_0 : boolean;
  signal type_cast_393_inst_req_1 : boolean;
  signal type_cast_331_inst_req_1 : boolean;
  signal addr_of_960_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_ack_0 : boolean;
  signal type_cast_1480_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_req_0 : boolean;
  signal type_cast_431_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_452_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_0 : boolean;
  signal type_cast_490_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 : boolean;
  signal addr_of_960_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1066_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_427_inst_ack_0 : boolean;
  signal type_cast_980_inst_req_1 : boolean;
  signal type_cast_980_inst_req_0 : boolean;
  signal type_cast_516_inst_req_0 : boolean;
  signal type_cast_516_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_ack_1 : boolean;
  signal type_cast_998_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_req_1 : boolean;
  signal type_cast_512_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_850_inst_req_0 : boolean;
  signal type_cast_481_inst_ack_1 : boolean;
  signal type_cast_551_inst_req_0 : boolean;
  signal type_cast_456_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal array_obj_ref_959_index_offset_req_1 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_req_1 : boolean;
  signal array_obj_ref_959_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_ack_1 : boolean;
  signal type_cast_512_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1084_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1030_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_427_inst_req_0 : boolean;
  signal type_cast_1034_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_439_inst_ack_0 : boolean;
  signal type_cast_456_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_ack_1 : boolean;
  signal type_cast_551_inst_req_1 : boolean;
  signal type_cast_836_inst_ack_1 : boolean;
  signal type_cast_490_inst_req_1 : boolean;
  signal type_cast_468_inst_ack_1 : boolean;
  signal type_cast_551_inst_ack_0 : boolean;
  signal type_cast_468_inst_req_1 : boolean;
  signal type_cast_1016_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1540_inst_req_0 : boolean;
  signal type_cast_494_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_464_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_1 : boolean;
  signal type_cast_538_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_439_inst_req_0 : boolean;
  signal type_cast_1070_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_464_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_ack_0 : boolean;
  signal type_cast_418_inst_ack_1 : boolean;
  signal type_cast_551_inst_ack_1 : boolean;
  signal type_cast_1034_inst_req_0 : boolean;
  signal type_cast_490_inst_ack_0 : boolean;
  signal type_cast_418_inst_req_1 : boolean;
  signal type_cast_343_inst_req_1 : boolean;
  signal type_cast_498_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_477_inst_ack_1 : boolean;
  signal type_cast_343_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_477_inst_req_1 : boolean;
  signal type_cast_498_inst_req_1 : boolean;
  signal type_cast_343_inst_req_0 : boolean;
  signal ptr_deref_880_store_0_ack_1 : boolean;
  signal type_cast_498_inst_ack_0 : boolean;
  signal type_cast_1500_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_ack_0 : boolean;
  signal type_cast_368_inst_ack_1 : boolean;
  signal type_cast_381_inst_ack_1 : boolean;
  signal type_cast_368_inst_req_1 : boolean;
  signal type_cast_368_inst_ack_0 : boolean;
  signal type_cast_368_inst_req_0 : boolean;
  signal type_cast_818_inst_req_0 : boolean;
  signal addr_of_960_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1048_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_314_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_314_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_314_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_314_inst_ack_1 : boolean;
  signal type_cast_318_inst_req_0 : boolean;
  signal type_cast_318_inst_ack_0 : boolean;
  signal type_cast_318_inst_req_1 : boolean;
  signal type_cast_318_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_327_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_327_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_327_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_327_inst_ack_1 : boolean;
  signal type_cast_836_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_559_inst_req_0 : boolean;
  signal array_obj_ref_959_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_559_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_559_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_559_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1084_inst_ack_0 : boolean;
  signal type_cast_1480_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1066_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1030_inst_ack_0 : boolean;
  signal type_cast_563_inst_req_0 : boolean;
  signal type_cast_563_inst_ack_0 : boolean;
  signal type_cast_563_inst_req_1 : boolean;
  signal type_cast_563_inst_ack_1 : boolean;
  signal type_cast_1088_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_ack_0 : boolean;
  signal type_cast_836_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1084_inst_req_0 : boolean;
  signal type_cast_1052_inst_ack_1 : boolean;
  signal type_cast_1052_inst_req_1 : boolean;
  signal type_cast_872_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1030_inst_req_0 : boolean;
  signal type_cast_576_inst_req_0 : boolean;
  signal type_cast_576_inst_ack_0 : boolean;
  signal type_cast_576_inst_req_1 : boolean;
  signal type_cast_576_inst_ack_1 : boolean;
  signal type_cast_1088_inst_req_0 : boolean;
  signal type_cast_836_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_584_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_584_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_584_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_584_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_976_inst_ack_1 : boolean;
  signal type_cast_872_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_976_inst_req_1 : boolean;
  signal type_cast_588_inst_req_0 : boolean;
  signal type_cast_588_inst_ack_0 : boolean;
  signal type_cast_588_inst_req_1 : boolean;
  signal type_cast_588_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_597_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_597_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_597_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_597_inst_ack_1 : boolean;
  signal type_cast_1052_inst_ack_0 : boolean;
  signal type_cast_1052_inst_req_0 : boolean;
  signal type_cast_872_inst_ack_0 : boolean;
  signal type_cast_872_inst_req_0 : boolean;
  signal type_cast_601_inst_req_0 : boolean;
  signal type_cast_601_inst_ack_0 : boolean;
  signal type_cast_601_inst_req_1 : boolean;
  signal type_cast_601_inst_ack_1 : boolean;
  signal type_cast_1399_inst_ack_1 : boolean;
  signal type_cast_1500_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_609_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_609_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_609_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_609_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1066_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_976_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_976_inst_req_0 : boolean;
  signal type_cast_613_inst_req_0 : boolean;
  signal type_cast_613_inst_ack_0 : boolean;
  signal type_cast_613_inst_req_1 : boolean;
  signal type_cast_613_inst_ack_1 : boolean;
  signal if_stmt_1377_branch_ack_0 : boolean;
  signal type_cast_1500_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_622_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_622_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_832_inst_ack_1 : boolean;
  signal type_cast_1034_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_622_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_622_inst_ack_1 : boolean;
  signal type_cast_1480_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1537_inst_req_0 : boolean;
  signal type_cast_626_inst_req_0 : boolean;
  signal type_cast_626_inst_ack_0 : boolean;
  signal type_cast_626_inst_req_1 : boolean;
  signal type_cast_626_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_832_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1367_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_994_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_634_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_634_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_634_inst_req_1 : boolean;
  signal type_cast_917_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_634_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1066_inst_req_0 : boolean;
  signal type_cast_638_inst_req_0 : boolean;
  signal type_cast_917_inst_req_1 : boolean;
  signal type_cast_638_inst_ack_0 : boolean;
  signal type_cast_638_inst_req_1 : boolean;
  signal type_cast_638_inst_ack_1 : boolean;
  signal type_cast_967_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_994_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_832_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_req_1 : boolean;
  signal type_cast_917_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_ack_1 : boolean;
  signal type_cast_1520_inst_req_0 : boolean;
  signal type_cast_967_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_868_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1361_inst_req_1 : boolean;
  signal type_cast_651_inst_req_0 : boolean;
  signal type_cast_917_inst_req_0 : boolean;
  signal type_cast_651_inst_ack_0 : boolean;
  signal type_cast_651_inst_req_1 : boolean;
  signal type_cast_651_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_832_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_868_inst_req_1 : boolean;
  signal type_cast_1070_inst_ack_1 : boolean;
  signal ptr_deref_880_store_0_ack_0 : boolean;
  signal if_stmt_664_branch_req_0 : boolean;
  signal ptr_deref_880_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_ack_1 : boolean;
  signal if_stmt_664_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_req_1 : boolean;
  signal if_stmt_664_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_850_inst_ack_1 : boolean;
  signal type_cast_967_inst_ack_0 : boolean;
  signal type_cast_1070_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1012_inst_ack_1 : boolean;
  signal if_stmt_679_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1531_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_ack_0 : boolean;
  signal if_stmt_679_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_req_0 : boolean;
  signal if_stmt_679_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_994_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_850_inst_req_1 : boolean;
  signal type_cast_967_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1012_inst_req_1 : boolean;
  signal type_cast_688_inst_req_0 : boolean;
  signal type_cast_688_inst_ack_0 : boolean;
  signal type_cast_688_inst_req_1 : boolean;
  signal type_cast_688_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_868_inst_ack_0 : boolean;
  signal type_cast_692_inst_req_0 : boolean;
  signal type_cast_692_inst_ack_0 : boolean;
  signal type_cast_1480_inst_req_1 : boolean;
  signal type_cast_692_inst_req_1 : boolean;
  signal type_cast_908_inst_ack_1 : boolean;
  signal type_cast_692_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_868_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1012_inst_ack_0 : boolean;
  signal type_cast_701_inst_req_0 : boolean;
  signal type_cast_908_inst_req_1 : boolean;
  signal type_cast_701_inst_ack_0 : boolean;
  signal type_cast_701_inst_req_1 : boolean;
  signal type_cast_701_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_994_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_963_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_963_inst_req_1 : boolean;
  signal array_obj_ref_743_index_offset_req_0 : boolean;
  signal array_obj_ref_743_index_offset_ack_0 : boolean;
  signal array_obj_ref_743_index_offset_req_1 : boolean;
  signal array_obj_ref_743_index_offset_ack_1 : boolean;
  signal type_cast_998_inst_ack_1 : boolean;
  signal type_cast_908_inst_ack_0 : boolean;
  signal type_cast_908_inst_req_0 : boolean;
  signal addr_of_744_final_reg_req_0 : boolean;
  signal addr_of_744_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1012_inst_req_0 : boolean;
  signal addr_of_744_final_reg_req_1 : boolean;
  signal addr_of_744_final_reg_ack_1 : boolean;
  signal type_cast_1070_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1531_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_963_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_963_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal type_cast_751_inst_req_1 : boolean;
  signal type_cast_751_inst_ack_1 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1048_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1048_inst_req_1 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1528_inst_req_1 : boolean;
  signal type_cast_764_inst_req_0 : boolean;
  signal if_stmt_894_branch_ack_0 : boolean;
  signal type_cast_764_inst_ack_0 : boolean;
  signal type_cast_764_inst_req_1 : boolean;
  signal type_cast_764_inst_ack_1 : boolean;
  signal type_cast_818_inst_ack_1 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 : boolean;
  signal type_cast_818_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_1 : boolean;
  signal if_stmt_894_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1048_inst_ack_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal type_cast_782_inst_req_0 : boolean;
  signal type_cast_782_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1528_inst_req_0 : boolean;
  signal type_cast_782_inst_req_1 : boolean;
  signal type_cast_782_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_0 : boolean;
  signal if_stmt_894_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 : boolean;
  signal type_cast_818_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1364_inst_ack_0 : boolean;
  signal type_cast_800_inst_req_0 : boolean;
  signal type_cast_800_inst_ack_0 : boolean;
  signal type_cast_1088_inst_req_1 : boolean;
  signal type_cast_1088_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1543_inst_ack_0 : boolean;
  signal type_cast_1470_inst_ack_1 : boolean;
  signal type_cast_1470_inst_req_1 : boolean;
  signal type_cast_1470_inst_ack_0 : boolean;
  signal if_stmt_1377_branch_ack_1 : boolean;
  signal type_cast_1399_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1367_inst_req_0 : boolean;
  signal type_cast_1490_inst_ack_1 : boolean;
  signal ptr_deref_1096_store_0_req_0 : boolean;
  signal ptr_deref_1096_store_0_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1361_inst_ack_0 : boolean;
  signal ptr_deref_1096_store_0_req_1 : boolean;
  signal ptr_deref_1096_store_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1543_inst_req_0 : boolean;
  signal if_stmt_1377_branch_req_0 : boolean;
  signal type_cast_1510_inst_ack_1 : boolean;
  signal type_cast_1490_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1361_inst_req_0 : boolean;
  signal if_stmt_1110_branch_req_0 : boolean;
  signal type_cast_1399_inst_ack_0 : boolean;
  signal if_stmt_1110_branch_ack_1 : boolean;
  signal type_cast_1399_inst_req_0 : boolean;
  signal if_stmt_1110_branch_ack_0 : boolean;
  signal type_cast_1510_inst_req_1 : boolean;
  signal type_cast_1470_inst_req_0 : boolean;
  signal type_cast_1121_inst_req_0 : boolean;
  signal type_cast_1121_inst_ack_0 : boolean;
  signal type_cast_1121_inst_req_1 : boolean;
  signal type_cast_1121_inst_ack_1 : boolean;
  signal type_cast_1125_inst_req_0 : boolean;
  signal type_cast_1125_inst_ack_0 : boolean;
  signal type_cast_1125_inst_req_1 : boolean;
  signal type_cast_1125_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1534_inst_ack_1 : boolean;
  signal type_cast_1129_inst_req_0 : boolean;
  signal type_cast_1129_inst_ack_0 : boolean;
  signal type_cast_1129_inst_req_1 : boolean;
  signal type_cast_1129_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1534_inst_req_1 : boolean;
  signal if_stmt_1147_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1373_inst_ack_1 : boolean;
  signal if_stmt_1147_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1358_inst_ack_1 : boolean;
  signal if_stmt_1147_branch_ack_0 : boolean;
  signal type_cast_1390_inst_ack_1 : boolean;
  signal type_cast_1156_inst_req_0 : boolean;
  signal type_cast_1156_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1525_inst_ack_1 : boolean;
  signal type_cast_1156_inst_req_1 : boolean;
  signal type_cast_1156_inst_ack_1 : boolean;
  signal type_cast_1460_inst_ack_1 : boolean;
  signal type_cast_1460_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1373_inst_req_1 : boolean;
  signal type_cast_1160_inst_req_0 : boolean;
  signal type_cast_1160_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1525_inst_req_1 : boolean;
  signal type_cast_1160_inst_req_1 : boolean;
  signal type_cast_1160_inst_ack_1 : boolean;
  signal type_cast_1169_inst_req_0 : boolean;
  signal type_cast_1169_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1525_inst_ack_0 : boolean;
  signal type_cast_1169_inst_req_1 : boolean;
  signal type_cast_1169_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1534_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1534_inst_req_0 : boolean;
  signal type_cast_1510_inst_ack_0 : boolean;
  signal type_cast_1510_inst_req_0 : boolean;
  signal type_cast_1460_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1373_inst_ack_0 : boolean;
  signal type_cast_1460_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1358_inst_req_1 : boolean;
  signal type_cast_1390_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1373_inst_req_0 : boolean;
  signal array_obj_ref_1211_index_offset_req_0 : boolean;
  signal array_obj_ref_1211_index_offset_ack_0 : boolean;
  signal array_obj_ref_1211_index_offset_req_1 : boolean;
  signal array_obj_ref_1211_index_offset_ack_1 : boolean;
  signal addr_of_1212_final_reg_req_0 : boolean;
  signal addr_of_1442_final_reg_ack_1 : boolean;
  signal addr_of_1212_final_reg_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1525_inst_req_0 : boolean;
  signal addr_of_1212_final_reg_req_1 : boolean;
  signal addr_of_1442_final_reg_req_1 : boolean;
  signal addr_of_1212_final_reg_ack_1 : boolean;
  signal type_cast_1450_inst_ack_1 : boolean;
  signal type_cast_1450_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1370_inst_ack_1 : boolean;
  signal addr_of_1442_final_reg_ack_0 : boolean;
  signal addr_of_1442_final_reg_req_0 : boolean;
  signal ptr_deref_1215_store_0_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1370_inst_req_1 : boolean;
  signal ptr_deref_1215_store_0_ack_0 : boolean;
  signal type_cast_1390_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1364_inst_ack_1 : boolean;
  signal ptr_deref_1215_store_0_req_1 : boolean;
  signal ptr_deref_1215_store_0_ack_1 : boolean;
  signal type_cast_1490_inst_ack_0 : boolean;
  signal type_cast_1390_inst_req_0 : boolean;
  signal if_stmt_1230_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1370_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1358_inst_ack_0 : boolean;
  signal if_stmt_1230_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1358_inst_req_0 : boolean;
  signal if_stmt_1230_branch_ack_0 : boolean;
  signal type_cast_1490_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1364_inst_req_1 : boolean;
  signal type_cast_1450_inst_ack_0 : boolean;
  signal call_stmt_1241_call_req_0 : boolean;
  signal call_stmt_1241_call_ack_0 : boolean;
  signal call_stmt_1241_call_req_1 : boolean;
  signal call_stmt_1241_call_ack_1 : boolean;
  signal type_cast_1450_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1370_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_req_1 : boolean;
  signal type_cast_1246_inst_req_0 : boolean;
  signal type_cast_1246_inst_ack_0 : boolean;
  signal type_cast_1246_inst_req_1 : boolean;
  signal type_cast_1246_inst_ack_1 : boolean;
  signal call_stmt_1263_call_req_0 : boolean;
  signal call_stmt_1263_call_ack_0 : boolean;
  signal type_cast_1386_inst_ack_1 : boolean;
  signal call_stmt_1263_call_req_1 : boolean;
  signal array_obj_ref_1441_index_offset_ack_1 : boolean;
  signal call_stmt_1263_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1540_inst_ack_1 : boolean;
  signal call_stmt_1266_call_req_0 : boolean;
  signal array_obj_ref_1441_index_offset_req_1 : boolean;
  signal call_stmt_1266_call_ack_0 : boolean;
  signal call_stmt_1266_call_req_1 : boolean;
  signal call_stmt_1266_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1540_inst_req_1 : boolean;
  signal type_cast_1386_inst_req_1 : boolean;
  signal type_cast_1270_inst_req_0 : boolean;
  signal array_obj_ref_1441_index_offset_ack_0 : boolean;
  signal type_cast_1270_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1522_inst_ack_1 : boolean;
  signal type_cast_1270_inst_req_1 : boolean;
  signal array_obj_ref_1441_index_offset_req_0 : boolean;
  signal type_cast_1270_inst_ack_1 : boolean;
  signal type_cast_1520_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1522_inst_req_1 : boolean;
  signal type_cast_1280_inst_req_0 : boolean;
  signal type_cast_1280_inst_ack_0 : boolean;
  signal type_cast_1280_inst_req_1 : boolean;
  signal type_cast_1280_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1537_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1528_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1522_inst_ack_0 : boolean;
  signal type_cast_1290_inst_req_0 : boolean;
  signal type_cast_1290_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1522_inst_req_0 : boolean;
  signal type_cast_1290_inst_req_1 : boolean;
  signal type_cast_1290_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1537_inst_req_1 : boolean;
  signal ptr_deref_1446_load_0_ack_1 : boolean;
  signal type_cast_1300_inst_req_0 : boolean;
  signal type_cast_1300_inst_ack_0 : boolean;
  signal type_cast_1300_inst_req_1 : boolean;
  signal type_cast_1300_inst_ack_1 : boolean;
  signal ptr_deref_1446_load_0_req_1 : boolean;
  signal type_cast_1310_inst_req_0 : boolean;
  signal type_cast_1310_inst_ack_0 : boolean;
  signal type_cast_1310_inst_req_1 : boolean;
  signal type_cast_1310_inst_ack_1 : boolean;
  signal type_cast_1320_inst_req_0 : boolean;
  signal type_cast_1320_inst_ack_0 : boolean;
  signal type_cast_1320_inst_req_1 : boolean;
  signal type_cast_1320_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1531_inst_ack_1 : boolean;
  signal ptr_deref_1446_load_0_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1367_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1540_inst_ack_0 : boolean;
  signal type_cast_1520_inst_ack_1 : boolean;
  signal type_cast_1330_inst_req_0 : boolean;
  signal type_cast_1330_inst_ack_0 : boolean;
  signal type_cast_1520_inst_req_1 : boolean;
  signal type_cast_1330_inst_req_1 : boolean;
  signal type_cast_1330_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1531_inst_req_1 : boolean;
  signal ptr_deref_1446_load_0_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1367_inst_req_1 : boolean;
  signal type_cast_1340_inst_req_0 : boolean;
  signal type_cast_1340_inst_ack_0 : boolean;
  signal type_cast_1340_inst_req_1 : boolean;
  signal type_cast_1340_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1537_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1361_inst_ack_1 : boolean;
  signal type_cast_1350_inst_req_0 : boolean;
  signal type_cast_1350_inst_ack_0 : boolean;
  signal type_cast_1350_inst_req_1 : boolean;
  signal type_cast_1350_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1352_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1355_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1543_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1543_inst_ack_1 : boolean;
  signal if_stmt_1557_branch_req_0 : boolean;
  signal if_stmt_1557_branch_ack_1 : boolean;
  signal if_stmt_1557_branch_ack_0 : boolean;
  signal phi_stmt_729_req_0 : boolean;
  signal type_cast_735_inst_req_0 : boolean;
  signal type_cast_735_inst_ack_0 : boolean;
  signal type_cast_735_inst_req_1 : boolean;
  signal type_cast_735_inst_ack_1 : boolean;
  signal phi_stmt_729_req_1 : boolean;
  signal phi_stmt_729_ack_0 : boolean;
  signal phi_stmt_945_req_1 : boolean;
  signal type_cast_948_inst_req_0 : boolean;
  signal type_cast_948_inst_ack_0 : boolean;
  signal type_cast_948_inst_req_1 : boolean;
  signal type_cast_948_inst_ack_1 : boolean;
  signal phi_stmt_945_req_0 : boolean;
  signal phi_stmt_945_ack_0 : boolean;
  signal phi_stmt_1197_req_0 : boolean;
  signal type_cast_1203_inst_req_0 : boolean;
  signal type_cast_1203_inst_ack_0 : boolean;
  signal type_cast_1203_inst_req_1 : boolean;
  signal type_cast_1203_inst_ack_1 : boolean;
  signal phi_stmt_1197_req_1 : boolean;
  signal phi_stmt_1197_ack_0 : boolean;
  signal phi_stmt_1427_req_0 : boolean;
  signal type_cast_1433_inst_req_0 : boolean;
  signal type_cast_1433_inst_ack_0 : boolean;
  signal type_cast_1433_inst_req_1 : boolean;
  signal type_cast_1433_inst_ack_1 : boolean;
  signal phi_stmt_1427_req_1 : boolean;
  signal phi_stmt_1427_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_772_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_772_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_772_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_772_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_772: Block -- control-path 
    signal convTranspose_CP_772_elements: BooleanArray(371 downto 0);
    -- 
  begin -- 
    convTranspose_CP_772_elements(0) <= convTranspose_CP_772_start;
    convTranspose_CP_772_symbol <= convTranspose_CP_772_elements(371);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	75 
    -- CP-element group 0: 	79 
    -- CP-element group 0: 	83 
    -- CP-element group 0: 	87 
    -- CP-element group 0: 	91 
    -- CP-element group 0: 	95 
    -- CP-element group 0: 	99 
    -- CP-element group 0: 	103 
    -- CP-element group 0: 	107 
    -- CP-element group 0: 	111 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0:  members (95) 
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_312/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/branch_block_stmt_312__entry__
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663__entry__
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_update_start_
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Update/cr
      -- 
    cr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_481_inst_req_1); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_431_inst_req_1); -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_356_inst_req_1); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_381_inst_req_1); -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_456_inst_req_1); -- 
    cr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_516_inst_req_1); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_443_inst_req_1); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_406_inst_req_1); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_393_inst_req_1); -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_331_inst_req_1); -- 
    cr_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_512_inst_req_1); -- 
    cr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_551_inst_req_1); -- 
    cr_1267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_490_inst_req_1); -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_468_inst_req_1); -- 
    cr_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_494_inst_req_1); -- 
    cr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_538_inst_req_1); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_418_inst_req_1); -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_343_inst_req_1); -- 
    cr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_498_inst_req_1); -- 
    cr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_368_inst_req_1); -- 
    rr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => RPIPE_ConvTranspose_input_pipe_314_inst_req_0); -- 
    cr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_318_inst_req_1); -- 
    cr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_563_inst_req_1); -- 
    cr_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_576_inst_req_1); -- 
    cr_1463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_588_inst_req_1); -- 
    cr_1491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_601_inst_req_1); -- 
    cr_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_613_inst_req_1); -- 
    cr_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_626_inst_req_1); -- 
    cr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_638_inst_req_1); -- 
    cr_1603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(0), ack => type_cast_651_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_update_start_
      -- CP-element group 1: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Update/cr
      -- 
    ra_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_314_inst_ack_0, ack => convTranspose_CP_772_elements(1)); -- 
    cr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(1), ack => RPIPE_ConvTranspose_input_pipe_314_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_314_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Sample/rr
      -- 
    ca_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_314_inst_ack_1, ack => convTranspose_CP_772_elements(2)); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(2), ack => type_cast_318_inst_req_0); -- 
    rr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(2), ack => RPIPE_ConvTranspose_input_pipe_327_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Sample/ra
      -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_318_inst_ack_0, ack => convTranspose_CP_772_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_318_Update/ca
      -- 
    ca_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_318_inst_ack_1, ack => convTranspose_CP_772_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_update_start_
      -- CP-element group 5: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Update/cr
      -- 
    ra_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_327_inst_ack_0, ack => convTranspose_CP_772_elements(5)); -- 
    cr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(5), ack => RPIPE_ConvTranspose_input_pipe_327_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_327_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Sample/$entry
      -- 
    ca_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_327_inst_ack_1, ack => convTranspose_CP_772_elements(6)); -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(6), ack => type_cast_331_inst_req_0); -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(6), ack => RPIPE_ConvTranspose_input_pipe_339_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_sample_completed_
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_331_inst_ack_0, ack => convTranspose_CP_772_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_331_update_completed_
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_331_inst_ack_1, ack => convTranspose_CP_772_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_update_start_
      -- CP-element group 9: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Sample/ra
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_339_inst_ack_0, ack => convTranspose_CP_772_elements(9)); -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(9), ack => RPIPE_ConvTranspose_input_pipe_339_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_339_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_sample_start_
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_339_inst_ack_1, ack => convTranspose_CP_772_elements(10)); -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(10), ack => type_cast_343_inst_req_0); -- 
    rr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(10), ack => RPIPE_ConvTranspose_input_pipe_352_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_sample_completed_
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_343_inst_ack_0, ack => convTranspose_CP_772_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_343_update_completed_
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_343_inst_ack_1, ack => convTranspose_CP_772_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_update_start_
      -- CP-element group 13: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Update/$entry
      -- 
    ra_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_352_inst_ack_0, ack => convTranspose_CP_772_elements(13)); -- 
    cr_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(13), ack => RPIPE_ConvTranspose_input_pipe_352_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_352_Update/$exit
      -- 
    ca_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_352_inst_ack_1, ack => convTranspose_CP_772_elements(14)); -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(14), ack => type_cast_356_inst_req_0); -- 
    rr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(14), ack => RPIPE_ConvTranspose_input_pipe_364_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_sample_completed_
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_356_inst_ack_0, ack => convTranspose_CP_772_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_356_Update/ca
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_356_inst_ack_1, ack => convTranspose_CP_772_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_update_start_
      -- CP-element group 17: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Sample/ra
      -- 
    ra_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_364_inst_ack_0, ack => convTranspose_CP_772_elements(17)); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(17), ack => RPIPE_ConvTranspose_input_pipe_364_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_364_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Sample/$entry
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_364_inst_ack_1, ack => convTranspose_CP_772_elements(18)); -- 
    rr_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(18), ack => type_cast_368_inst_req_0); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(18), ack => RPIPE_ConvTranspose_input_pipe_377_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Sample/$exit
      -- 
    ra_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_0, ack => convTranspose_CP_772_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_368_update_completed_
      -- 
    ca_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_1, ack => convTranspose_CP_772_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_update_start_
      -- CP-element group 21: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_sample_completed_
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_377_inst_ack_0, ack => convTranspose_CP_772_elements(21)); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(21), ack => RPIPE_ConvTranspose_input_pipe_377_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_377_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_sample_start_
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_377_inst_ack_1, ack => convTranspose_CP_772_elements(22)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(22), ack => type_cast_381_inst_req_0); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(22), ack => RPIPE_ConvTranspose_input_pipe_389_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_sample_completed_
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_381_inst_ack_0, ack => convTranspose_CP_772_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_381_Update/ca
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_381_inst_ack_1, ack => convTranspose_CP_772_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_update_start_
      -- CP-element group 25: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_sample_completed_
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_389_inst_ack_0, ack => convTranspose_CP_772_elements(25)); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(25), ack => RPIPE_ConvTranspose_input_pipe_389_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_389_update_completed_
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_389_inst_ack_1, ack => convTranspose_CP_772_elements(26)); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(26), ack => RPIPE_ConvTranspose_input_pipe_402_inst_req_0); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(26), ack => type_cast_393_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Sample/$exit
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_393_inst_ack_0, ack => convTranspose_CP_772_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	112 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_393_Update/$exit
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_393_inst_ack_1, ack => convTranspose_CP_772_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_update_start_
      -- CP-element group 29: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Update/cr
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_402_inst_ack_0, ack => convTranspose_CP_772_elements(29)); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(29), ack => RPIPE_ConvTranspose_input_pipe_402_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_402_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_sample_start_
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_402_inst_ack_1, ack => convTranspose_CP_772_elements(30)); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(30), ack => RPIPE_ConvTranspose_input_pipe_414_inst_req_0); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(30), ack => type_cast_406_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_sample_completed_
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_406_inst_ack_0, ack => convTranspose_CP_772_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	112 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_406_Update/$exit
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_406_inst_ack_1, ack => convTranspose_CP_772_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_update_start_
      -- CP-element group 33: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Sample/ra
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_414_inst_ack_0, ack => convTranspose_CP_772_elements(33)); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(33), ack => RPIPE_ConvTranspose_input_pipe_414_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_414_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_sample_start_
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_414_inst_ack_1, ack => convTranspose_CP_772_elements(34)); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(34), ack => RPIPE_ConvTranspose_input_pipe_427_inst_req_0); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(34), ack => type_cast_418_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Sample/ra
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_418_inst_ack_0, ack => convTranspose_CP_772_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	66 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_418_Update/ca
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_418_inst_ack_1, ack => convTranspose_CP_772_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_update_start_
      -- CP-element group 37: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_sample_completed_
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_427_inst_ack_0, ack => convTranspose_CP_772_elements(37)); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(37), ack => RPIPE_ConvTranspose_input_pipe_427_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_427_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Sample/rr
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_427_inst_ack_1, ack => convTranspose_CP_772_elements(38)); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(38), ack => type_cast_431_inst_req_0); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(38), ack => RPIPE_ConvTranspose_input_pipe_439_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Sample/ra
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_431_inst_ack_0, ack => convTranspose_CP_772_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	66 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_431_Update/ca
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_431_inst_ack_1, ack => convTranspose_CP_772_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_update_start_
      -- CP-element group 41: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Sample/ra
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_439_inst_ack_0, ack => convTranspose_CP_772_elements(41)); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(41), ack => RPIPE_ConvTranspose_input_pipe_439_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_439_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Sample/$entry
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_439_inst_ack_1, ack => convTranspose_CP_772_elements(42)); -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(42), ack => type_cast_443_inst_req_0); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(42), ack => RPIPE_ConvTranspose_input_pipe_452_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Sample/$exit
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_0, ack => convTranspose_CP_772_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	69 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_443_update_completed_
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_1, ack => convTranspose_CP_772_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_update_start_
      -- CP-element group 45: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Update/cr
      -- CP-element group 45: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_sample_completed_
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_452_inst_ack_0, ack => convTranspose_CP_772_elements(45)); -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(45), ack => RPIPE_ConvTranspose_input_pipe_452_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_452_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Sample/rr
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_452_inst_ack_1, ack => convTranspose_CP_772_elements(46)); -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(46), ack => RPIPE_ConvTranspose_input_pipe_464_inst_req_0); -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(46), ack => type_cast_456_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Sample/$exit
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_0, ack => convTranspose_CP_772_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	69 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_456_update_completed_
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_1, ack => convTranspose_CP_772_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_update_start_
      -- CP-element group 49: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Sample/$exit
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_464_inst_ack_0, ack => convTranspose_CP_772_elements(49)); -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(49), ack => RPIPE_ConvTranspose_input_pipe_464_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_464_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Sample/$entry
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_464_inst_ack_1, ack => convTranspose_CP_772_elements(50)); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(50), ack => type_cast_468_inst_req_0); -- 
    rr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(50), ack => RPIPE_ConvTranspose_input_pipe_477_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Sample/$exit
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_468_inst_ack_0, ack => convTranspose_CP_772_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	112 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_468_Update/$exit
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_468_inst_ack_1, ack => convTranspose_CP_772_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_update_start_
      -- CP-element group 53: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Update/$entry
      -- 
    ra_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_477_inst_ack_0, ack => convTranspose_CP_772_elements(53)); -- 
    cr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(53), ack => RPIPE_ConvTranspose_input_pipe_477_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	72 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_477_Update/$exit
      -- 
    ca_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_477_inst_ack_1, ack => convTranspose_CP_772_elements(54)); -- 
    rr_1248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(54), ack => type_cast_481_inst_req_0); -- 
    rr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(54), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Sample/$exit
      -- 
    ra_1249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_0, ack => convTranspose_CP_772_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	112 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_481_Update/ca
      -- 
    ca_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_1, ack => convTranspose_CP_772_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Sample/$entry
      -- 
    rr_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(57), ack => type_cast_490_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(4) & convTranspose_CP_772_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Sample/ra
      -- 
    ra_1263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_0, ack => convTranspose_CP_772_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	112 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_490_update_completed_
      -- 
    ca_1268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_1, ack => convTranspose_CP_772_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Sample/$entry
      -- 
    rr_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(60), ack => type_cast_494_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(12) & convTranspose_CP_772_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Sample/ra
      -- 
    ra_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_0, ack => convTranspose_CP_772_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	112 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_494_update_completed_
      -- 
    ca_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_1, ack => convTranspose_CP_772_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Sample/$entry
      -- 
    rr_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(63), ack => type_cast_498_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(20) & convTranspose_CP_772_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Sample/ra
      -- 
    ra_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_0, ack => convTranspose_CP_772_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	112 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_498_Update/ca
      -- 
    ca_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_1, ack => convTranspose_CP_772_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	36 
    -- CP-element group 66: 	40 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_sample_start_
      -- 
    rr_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(66), ack => type_cast_512_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(36) & convTranspose_CP_772_elements(40);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_sample_completed_
      -- 
    ra_1305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_512_inst_ack_0, ack => convTranspose_CP_772_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	112 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_512_update_completed_
      -- 
    ca_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_512_inst_ack_1, ack => convTranspose_CP_772_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	44 
    -- CP-element group 69: 	48 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Sample/$entry
      -- 
    rr_1318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(69), ack => type_cast_516_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(44) & convTranspose_CP_772_elements(48);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_sample_completed_
      -- 
    ra_1319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_516_inst_ack_0, ack => convTranspose_CP_772_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	112 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_516_update_completed_
      -- 
    ca_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_516_inst_ack_1, ack => convTranspose_CP_772_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	54 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_update_start_
      -- 
    ra_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_0, ack => convTranspose_CP_772_elements(72)); -- 
    cr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(72), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_1); -- 
    -- CP-element group 73:  fork  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	76 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_534_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Sample/rr
      -- 
    ca_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_1, ack => convTranspose_CP_772_elements(73)); -- 
    rr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(73), ack => type_cast_538_inst_req_0); -- 
    rr_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(73), ack => RPIPE_ConvTranspose_input_pipe_547_inst_req_0); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Sample/$exit
      -- 
    ra_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => convTranspose_CP_772_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	0 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	112 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_538_update_completed_
      -- 
    ca_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_1, ack => convTranspose_CP_772_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	73 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_update_start_
      -- CP-element group 76: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_sample_completed_
      -- 
    ra_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_547_inst_ack_0, ack => convTranspose_CP_772_elements(76)); -- 
    cr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(76), ack => RPIPE_ConvTranspose_input_pipe_547_inst_req_1); -- 
    -- CP-element group 77:  fork  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	80 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_547_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Sample/rr
      -- 
    ca_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_547_inst_ack_1, ack => convTranspose_CP_772_elements(77)); -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(77), ack => type_cast_551_inst_req_0); -- 
    rr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(77), ack => RPIPE_ConvTranspose_input_pipe_559_inst_req_0); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_sample_completed_
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_551_inst_ack_0, ack => convTranspose_CP_772_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	0 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	112 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_551_update_completed_
      -- 
    ca_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_551_inst_ack_1, ack => convTranspose_CP_772_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	77 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_update_start_
      -- CP-element group 80: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Update/cr
      -- 
    ra_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_559_inst_ack_0, ack => convTranspose_CP_772_elements(80)); -- 
    cr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(80), ack => RPIPE_ConvTranspose_input_pipe_559_inst_req_1); -- 
    -- CP-element group 81:  fork  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: 	84 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_559_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Sample/rr
      -- 
    ca_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_559_inst_ack_1, ack => convTranspose_CP_772_elements(81)); -- 
    rr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(81), ack => type_cast_563_inst_req_0); -- 
    rr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(81), ack => RPIPE_ConvTranspose_input_pipe_572_inst_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Sample/ra
      -- 
    ra_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_563_inst_ack_0, ack => convTranspose_CP_772_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	0 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	112 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_563_Update/ca
      -- 
    ca_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_563_inst_ack_1, ack => convTranspose_CP_772_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	81 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_update_start_
      -- CP-element group 84: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Update/cr
      -- 
    ra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_572_inst_ack_0, ack => convTranspose_CP_772_elements(84)); -- 
    cr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(84), ack => RPIPE_ConvTranspose_input_pipe_572_inst_req_1); -- 
    -- CP-element group 85:  fork  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	88 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_572_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Sample/rr
      -- 
    ca_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_572_inst_ack_1, ack => convTranspose_CP_772_elements(85)); -- 
    rr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(85), ack => type_cast_576_inst_req_0); -- 
    rr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(85), ack => RPIPE_ConvTranspose_input_pipe_584_inst_req_0); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Sample/ra
      -- 
    ra_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_576_inst_ack_0, ack => convTranspose_CP_772_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	0 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	112 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_576_Update/ca
      -- 
    ca_1436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_576_inst_ack_1, ack => convTranspose_CP_772_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	85 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_update_start_
      -- CP-element group 88: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Update/cr
      -- 
    ra_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_584_inst_ack_0, ack => convTranspose_CP_772_elements(88)); -- 
    cr_1449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(88), ack => RPIPE_ConvTranspose_input_pipe_584_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (9) 
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_584_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Sample/rr
      -- 
    ca_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_584_inst_ack_1, ack => convTranspose_CP_772_elements(89)); -- 
    rr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(89), ack => type_cast_588_inst_req_0); -- 
    rr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(89), ack => RPIPE_ConvTranspose_input_pipe_597_inst_req_0); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Sample/ra
      -- 
    ra_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_588_inst_ack_0, ack => convTranspose_CP_772_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	0 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	112 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_588_Update/ca
      -- 
    ca_1464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_588_inst_ack_1, ack => convTranspose_CP_772_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	89 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_update_start_
      -- CP-element group 92: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Update/cr
      -- 
    ra_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_597_inst_ack_0, ack => convTranspose_CP_772_elements(92)); -- 
    cr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(92), ack => RPIPE_ConvTranspose_input_pipe_597_inst_req_1); -- 
    -- CP-element group 93:  fork  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: 	96 
    -- CP-element group 93:  members (9) 
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_597_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Sample/rr
      -- 
    ca_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_597_inst_ack_1, ack => convTranspose_CP_772_elements(93)); -- 
    rr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(93), ack => type_cast_601_inst_req_0); -- 
    rr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(93), ack => RPIPE_ConvTranspose_input_pipe_609_inst_req_0); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Sample/ra
      -- 
    ra_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_0, ack => convTranspose_CP_772_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	0 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	112 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_601_Update/ca
      -- 
    ca_1492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_1, ack => convTranspose_CP_772_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	93 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_update_start_
      -- CP-element group 96: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Update/cr
      -- 
    ra_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_609_inst_ack_0, ack => convTranspose_CP_772_elements(96)); -- 
    cr_1505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(96), ack => RPIPE_ConvTranspose_input_pipe_609_inst_req_1); -- 
    -- CP-element group 97:  fork  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (9) 
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_609_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Sample/rr
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Sample/rr
      -- 
    ca_1506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_609_inst_ack_1, ack => convTranspose_CP_772_elements(97)); -- 
    rr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(97), ack => type_cast_613_inst_req_0); -- 
    rr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(97), ack => RPIPE_ConvTranspose_input_pipe_622_inst_req_0); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Sample/ra
      -- 
    ra_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_0, ack => convTranspose_CP_772_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	0 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	112 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_613_Update/ca
      -- 
    ca_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_1, ack => convTranspose_CP_772_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_update_start_
      -- CP-element group 100: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Update/cr
      -- 
    ra_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_622_inst_ack_0, ack => convTranspose_CP_772_elements(100)); -- 
    cr_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(100), ack => RPIPE_ConvTranspose_input_pipe_622_inst_req_1); -- 
    -- CP-element group 101:  fork  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (9) 
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_622_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Sample/rr
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Sample/rr
      -- 
    ca_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_622_inst_ack_1, ack => convTranspose_CP_772_elements(101)); -- 
    rr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(101), ack => type_cast_626_inst_req_0); -- 
    rr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(101), ack => RPIPE_ConvTranspose_input_pipe_634_inst_req_0); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Sample/ra
      -- 
    ra_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_0, ack => convTranspose_CP_772_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	0 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	112 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_626_Update/ca
      -- 
    ca_1548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_1, ack => convTranspose_CP_772_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	101 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_update_start_
      -- CP-element group 104: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Update/cr
      -- 
    ra_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_634_inst_ack_0, ack => convTranspose_CP_772_elements(104)); -- 
    cr_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(104), ack => RPIPE_ConvTranspose_input_pipe_634_inst_req_1); -- 
    -- CP-element group 105:  fork  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (9) 
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_634_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Sample/rr
      -- 
    ca_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_634_inst_ack_1, ack => convTranspose_CP_772_elements(105)); -- 
    rr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(105), ack => type_cast_638_inst_req_0); -- 
    rr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(105), ack => RPIPE_ConvTranspose_input_pipe_647_inst_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Sample/ra
      -- 
    ra_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_638_inst_ack_0, ack => convTranspose_CP_772_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	0 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_638_Update/ca
      -- 
    ca_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_638_inst_ack_1, ack => convTranspose_CP_772_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (6) 
      -- CP-element group 108: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_update_start_
      -- CP-element group 108: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Update/cr
      -- 
    ra_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_647_inst_ack_0, ack => convTranspose_CP_772_elements(108)); -- 
    cr_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(108), ack => RPIPE_ConvTranspose_input_pipe_647_inst_req_1); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/RPIPE_ConvTranspose_input_pipe_647_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Sample/rr
      -- 
    ca_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_647_inst_ack_1, ack => convTranspose_CP_772_elements(109)); -- 
    rr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(109), ack => type_cast_651_inst_req_0); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Sample/ra
      -- 
    ra_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_651_inst_ack_0, ack => convTranspose_CP_772_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	0 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/type_cast_651_Update/ca
      -- 
    ca_1604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_651_inst_ack_1, ack => convTranspose_CP_772_elements(111)); -- 
    -- CP-element group 112:  branch  join  transition  place  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	32 
    -- CP-element group 112: 	28 
    -- CP-element group 112: 	56 
    -- CP-element group 112: 	62 
    -- CP-element group 112: 	59 
    -- CP-element group 112: 	65 
    -- CP-element group 112: 	52 
    -- CP-element group 112: 	68 
    -- CP-element group 112: 	71 
    -- CP-element group 112: 	75 
    -- CP-element group 112: 	79 
    -- CP-element group 112: 	83 
    -- CP-element group 112: 	87 
    -- CP-element group 112: 	91 
    -- CP-element group 112: 	95 
    -- CP-element group 112: 	99 
    -- CP-element group 112: 	103 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (10) 
      -- CP-element group 112: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663__exit__
      -- CP-element group 112: 	 branch_block_stmt_312/if_stmt_664__entry__
      -- CP-element group 112: 	 branch_block_stmt_312/assign_stmt_315_to_assign_stmt_663/$exit
      -- CP-element group 112: 	 branch_block_stmt_312/if_stmt_664_dead_link/$entry
      -- CP-element group 112: 	 branch_block_stmt_312/if_stmt_664_eval_test/$entry
      -- CP-element group 112: 	 branch_block_stmt_312/if_stmt_664_eval_test/$exit
      -- CP-element group 112: 	 branch_block_stmt_312/if_stmt_664_eval_test/branch_req
      -- CP-element group 112: 	 branch_block_stmt_312/R_cmp430_665_place
      -- CP-element group 112: 	 branch_block_stmt_312/if_stmt_664_if_link/$entry
      -- CP-element group 112: 	 branch_block_stmt_312/if_stmt_664_else_link/$entry
      -- 
    branch_req_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(112), ack => if_stmt_664_branch_req_0); -- 
    convTranspose_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 18) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1);
      constant place_markings: IntegerArray(0 to 18)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0);
      constant place_delays: IntegerArray(0 to 18) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 19); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(32) & convTranspose_CP_772_elements(28) & convTranspose_CP_772_elements(56) & convTranspose_CP_772_elements(62) & convTranspose_CP_772_elements(59) & convTranspose_CP_772_elements(65) & convTranspose_CP_772_elements(52) & convTranspose_CP_772_elements(68) & convTranspose_CP_772_elements(71) & convTranspose_CP_772_elements(75) & convTranspose_CP_772_elements(79) & convTranspose_CP_772_elements(83) & convTranspose_CP_772_elements(87) & convTranspose_CP_772_elements(91) & convTranspose_CP_772_elements(95) & convTranspose_CP_772_elements(99) & convTranspose_CP_772_elements(103) & convTranspose_CP_772_elements(107) & convTranspose_CP_772_elements(111);
      gj_convTranspose_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 19, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	117 
    -- CP-element group 113: 	118 
    -- CP-element group 113: 	119 
    -- CP-element group 113: 	120 
    -- CP-element group 113: 	121 
    -- CP-element group 113: 	122 
    -- CP-element group 113:  members (30) 
      -- CP-element group 113: 	 branch_block_stmt_312/merge_stmt_685__exit__
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726__entry__
      -- CP-element group 113: 	 branch_block_stmt_312/if_stmt_664_if_link/$exit
      -- CP-element group 113: 	 branch_block_stmt_312/if_stmt_664_if_link/if_choice_transition
      -- CP-element group 113: 	 branch_block_stmt_312/entry_bbx_xnph432
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_update_start_
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_update_start_
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_update_start_
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_312/entry_bbx_xnph432_PhiReq/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/entry_bbx_xnph432_PhiReq/$exit
      -- CP-element group 113: 	 branch_block_stmt_312/merge_stmt_685_PhiReqMerge
      -- CP-element group 113: 	 branch_block_stmt_312/merge_stmt_685_PhiAck/$entry
      -- CP-element group 113: 	 branch_block_stmt_312/merge_stmt_685_PhiAck/$exit
      -- CP-element group 113: 	 branch_block_stmt_312/merge_stmt_685_PhiAck/dummy
      -- 
    if_choice_transition_1617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_664_branch_ack_1, ack => convTranspose_CP_772_elements(113)); -- 
    rr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(113), ack => type_cast_688_inst_req_0); -- 
    cr_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(113), ack => type_cast_688_inst_req_1); -- 
    rr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(113), ack => type_cast_692_inst_req_0); -- 
    cr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(113), ack => type_cast_692_inst_req_1); -- 
    rr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(113), ack => type_cast_701_inst_req_0); -- 
    cr_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(113), ack => type_cast_701_inst_req_1); -- 
    -- CP-element group 114:  transition  place  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	344 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_312/if_stmt_664_else_link/$exit
      -- CP-element group 114: 	 branch_block_stmt_312/if_stmt_664_else_link/else_choice_transition
      -- CP-element group 114: 	 branch_block_stmt_312/entry_forx_xcond176x_xpreheader
      -- CP-element group 114: 	 branch_block_stmt_312/entry_forx_xcond176x_xpreheader_PhiReq/$entry
      -- CP-element group 114: 	 branch_block_stmt_312/entry_forx_xcond176x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_1621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_664_branch_ack_0, ack => convTranspose_CP_772_elements(114)); -- 
    -- CP-element group 115:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	344 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	166 
    -- CP-element group 115: 	167 
    -- CP-element group 115: 	168 
    -- CP-element group 115: 	169 
    -- CP-element group 115:  members (24) 
      -- CP-element group 115: 	 branch_block_stmt_312/merge_stmt_900__exit__
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942__entry__
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_312/if_stmt_679_if_link/$exit
      -- CP-element group 115: 	 branch_block_stmt_312/if_stmt_679_if_link/if_choice_transition
      -- CP-element group 115: 	 branch_block_stmt_312/forx_xcond176x_xpreheader_bbx_xnph428
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_update_start_
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_update_start_
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/$entry
      -- CP-element group 115: 	 branch_block_stmt_312/forx_xcond176x_xpreheader_bbx_xnph428_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_312/forx_xcond176x_xpreheader_bbx_xnph428_PhiReq/$exit
      -- CP-element group 115: 	 branch_block_stmt_312/merge_stmt_900_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_312/merge_stmt_900_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_312/merge_stmt_900_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_312/merge_stmt_900_PhiAck/dummy
      -- 
    if_choice_transition_1639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_679_branch_ack_1, ack => convTranspose_CP_772_elements(115)); -- 
    cr_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(115), ack => type_cast_917_inst_req_1); -- 
    rr_2057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(115), ack => type_cast_917_inst_req_0); -- 
    cr_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(115), ack => type_cast_908_inst_req_1); -- 
    rr_2043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(115), ack => type_cast_908_inst_req_0); -- 
    -- CP-element group 116:  transition  place  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	344 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	357 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_312/if_stmt_679_else_link/$exit
      -- CP-element group 116: 	 branch_block_stmt_312/if_stmt_679_else_link/else_choice_transition
      -- CP-element group 116: 	 branch_block_stmt_312/forx_xcond176x_xpreheader_forx_xend235
      -- CP-element group 116: 	 branch_block_stmt_312/forx_xcond176x_xpreheader_forx_xend235_PhiReq/$entry
      -- CP-element group 116: 	 branch_block_stmt_312/forx_xcond176x_xpreheader_forx_xend235_PhiReq/$exit
      -- 
    else_choice_transition_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_679_branch_ack_0, ack => convTranspose_CP_772_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	113 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Sample/ra
      -- 
    ra_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_0, ack => convTranspose_CP_772_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	113 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_688_Update/ca
      -- 
    ca_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_1, ack => convTranspose_CP_772_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	113 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Sample/ra
      -- 
    ra_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_692_inst_ack_0, ack => convTranspose_CP_772_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_692_Update/ca
      -- 
    ca_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_692_inst_ack_1, ack => convTranspose_CP_772_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	113 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Sample/ra
      -- 
    ra_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_0, ack => convTranspose_CP_772_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	113 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/type_cast_701_Update/ca
      -- 
    ca_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_1, ack => convTranspose_CP_772_elements(122)); -- 
    -- CP-element group 123:  join  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	345 
    -- CP-element group 123:  members (6) 
      -- CP-element group 123: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726__exit__
      -- CP-element group 123: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody
      -- CP-element group 123: 	 branch_block_stmt_312/assign_stmt_689_to_assign_stmt_726/$exit
      -- CP-element group 123: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/phi_stmt_729/$entry
      -- CP-element group 123: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/$entry
      -- 
    convTranspose_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(118) & convTranspose_CP_772_elements(120) & convTranspose_CP_772_elements(122);
      gj_convTranspose_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	350 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	163 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_sample_complete
      -- CP-element group 124: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Sample/ack
      -- 
    ack_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_743_index_offset_ack_0, ack => convTranspose_CP_772_elements(124)); -- 
    -- CP-element group 125:  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	350 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (11) 
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_root_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_offset_calculated
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Update/ack
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_base_plus_offset/$entry
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_base_plus_offset/$exit
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_base_plus_offset/sum_rename_req
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_base_plus_offset/sum_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_request/$entry
      -- CP-element group 125: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_request/req
      -- 
    ack_1724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_743_index_offset_ack_1, ack => convTranspose_CP_772_elements(125)); -- 
    req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(125), ack => addr_of_744_final_reg_req_0); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_request/$exit
      -- CP-element group 126: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_request/ack
      -- 
    ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_744_final_reg_ack_0, ack => convTranspose_CP_772_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	350 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	160 
    -- CP-element group 127:  members (19) 
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_plus_offset/sum_rename_ack
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_plus_offset/sum_rename_req
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_addr_resize/base_resize_req
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_plus_offset/$exit
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_word_addrgen/$entry
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_plus_offset/$entry
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_addr_resize/$exit
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_word_addrgen/$exit
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_addr_resize/base_resize_ack
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_word_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_addr_resize/$entry
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_base_address_resized
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_root_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_word_addrgen/root_register_req
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_word_addrgen/root_register_ack
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_complete/$exit
      -- CP-element group 127: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_complete/ack
      -- 
    ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_744_final_reg_ack_1, ack => convTranspose_CP_772_elements(127)); -- 
    -- CP-element group 128:  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	350 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_update_start_
      -- CP-element group 128: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Sample/ra
      -- CP-element group 128: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Update/cr
      -- 
    ra_1748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_747_inst_ack_0, ack => convTranspose_CP_772_elements(128)); -- 
    cr_1752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(128), ack => RPIPE_ConvTranspose_input_pipe_747_inst_req_1); -- 
    -- CP-element group 129:  fork  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: 	132 
    -- CP-element group 129:  members (9) 
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Update/ca
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Sample/rr
      -- 
    ca_1753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_747_inst_ack_1, ack => convTranspose_CP_772_elements(129)); -- 
    rr_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(129), ack => type_cast_751_inst_req_0); -- 
    rr_1775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(129), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_0); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Sample/ra
      -- 
    ra_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => convTranspose_CP_772_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	350 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	160 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Update/ca
      -- 
    ca_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_1, ack => convTranspose_CP_772_elements(131)); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	129 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_update_start_
      -- CP-element group 132: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Sample/ra
      -- CP-element group 132: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Update/cr
      -- 
    ra_1776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_0, ack => convTranspose_CP_772_elements(132)); -- 
    cr_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(132), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_1); -- 
    -- CP-element group 133:  fork  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133: 	136 
    -- CP-element group 133:  members (9) 
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_760_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Sample/rr
      -- 
    ca_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_1, ack => convTranspose_CP_772_elements(133)); -- 
    rr_1789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(133), ack => type_cast_764_inst_req_0); -- 
    rr_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(133), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_0); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Sample/ra
      -- 
    ra_1790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_0, ack => convTranspose_CP_772_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	350 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	160 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Update/ca
      -- 
    ca_1795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_1, ack => convTranspose_CP_772_elements(135)); -- 
    -- CP-element group 136:  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	133 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (6) 
      -- CP-element group 136: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_update_start_
      -- CP-element group 136: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Sample/ra
      -- CP-element group 136: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Update/cr
      -- 
    ra_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_0, ack => convTranspose_CP_772_elements(136)); -- 
    cr_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(136), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_1); -- 
    -- CP-element group 137:  fork  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	140 
    -- CP-element group 137:  members (9) 
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_778_Update/ca
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Sample/rr
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Sample/rr
      -- 
    ca_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_1, ack => convTranspose_CP_772_elements(137)); -- 
    rr_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(137), ack => type_cast_782_inst_req_0); -- 
    rr_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(137), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_0); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Sample/ra
      -- 
    ra_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_0, ack => convTranspose_CP_772_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	350 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	160 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Update/ca
      -- 
    ca_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_1, ack => convTranspose_CP_772_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	137 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (6) 
      -- CP-element group 140: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_update_start_
      -- CP-element group 140: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Sample/ra
      -- CP-element group 140: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Update/cr
      -- 
    ra_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_0, ack => convTranspose_CP_772_elements(140)); -- 
    cr_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(140), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_1); -- 
    -- CP-element group 141:  fork  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141: 	144 
    -- CP-element group 141:  members (9) 
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_796_Update/ca
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Sample/rr
      -- 
    ca_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_1, ack => convTranspose_CP_772_elements(141)); -- 
    rr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(141), ack => type_cast_800_inst_req_0); -- 
    rr_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(141), ack => RPIPE_ConvTranspose_input_pipe_814_inst_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Sample/ra
      -- 
    ra_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_0, ack => convTranspose_CP_772_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	350 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	160 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_update_completed_
      -- 
    ca_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_1, ack => convTranspose_CP_772_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	141 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_update_start_
      -- CP-element group 144: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Sample/ra
      -- CP-element group 144: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Sample/$exit
      -- 
    ra_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_814_inst_ack_0, ack => convTranspose_CP_772_elements(144)); -- 
    cr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(144), ack => RPIPE_ConvTranspose_input_pipe_814_inst_req_1); -- 
    -- CP-element group 145:  fork  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145: 	148 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Update/ca
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_814_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_sample_start_
      -- 
    ca_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_814_inst_ack_1, ack => convTranspose_CP_772_elements(145)); -- 
    rr_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(145), ack => type_cast_818_inst_req_0); -- 
    rr_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(145), ack => RPIPE_ConvTranspose_input_pipe_832_inst_req_0); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Sample/ra
      -- 
    ra_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_0, ack => convTranspose_CP_772_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	350 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	160 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Update/$exit
      -- 
    ca_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_1, ack => convTranspose_CP_772_elements(147)); -- 
    -- CP-element group 148:  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	145 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Update/cr
      -- CP-element group 148: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Sample/ra
      -- CP-element group 148: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_update_start_
      -- CP-element group 148: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_sample_completed_
      -- 
    ra_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_832_inst_ack_0, ack => convTranspose_CP_772_elements(148)); -- 
    cr_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(148), ack => RPIPE_ConvTranspose_input_pipe_832_inst_req_1); -- 
    -- CP-element group 149:  fork  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	152 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Update/ca
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_832_update_completed_
      -- 
    ca_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_832_inst_ack_1, ack => convTranspose_CP_772_elements(149)); -- 
    rr_1901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(149), ack => type_cast_836_inst_req_0); -- 
    rr_1915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(149), ack => RPIPE_ConvTranspose_input_pipe_850_inst_req_0); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_sample_completed_
      -- 
    ra_1902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_836_inst_ack_0, ack => convTranspose_CP_772_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	350 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	160 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_update_completed_
      -- 
    ca_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_836_inst_ack_1, ack => convTranspose_CP_772_elements(151)); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	149 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_update_start_
      -- CP-element group 152: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Update/cr
      -- 
    ra_1916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_850_inst_ack_0, ack => convTranspose_CP_772_elements(152)); -- 
    cr_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(152), ack => RPIPE_ConvTranspose_input_pipe_850_inst_req_1); -- 
    -- CP-element group 153:  fork  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	156 
    -- CP-element group 153:  members (9) 
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_850_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Sample/$entry
      -- 
    ca_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_850_inst_ack_1, ack => convTranspose_CP_772_elements(153)); -- 
    rr_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(153), ack => type_cast_854_inst_req_0); -- 
    rr_1943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(153), ack => RPIPE_ConvTranspose_input_pipe_868_inst_req_0); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Sample/$exit
      -- 
    ra_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => convTranspose_CP_772_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	350 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	160 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_update_completed_
      -- 
    ca_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => convTranspose_CP_772_elements(155)); -- 
    -- CP-element group 156:  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (6) 
      -- CP-element group 156: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_update_start_
      -- CP-element group 156: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_sample_completed_
      -- 
    ra_1944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_868_inst_ack_0, ack => convTranspose_CP_772_elements(156)); -- 
    cr_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(156), ack => RPIPE_ConvTranspose_input_pipe_868_inst_req_1); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Sample/rr
      -- CP-element group 157: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_868_update_completed_
      -- 
    ca_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_868_inst_ack_1, ack => convTranspose_CP_772_elements(157)); -- 
    rr_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(157), ack => type_cast_872_inst_req_0); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_sample_completed_
      -- 
    ra_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_872_inst_ack_0, ack => convTranspose_CP_772_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	350 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_update_completed_
      -- 
    ca_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_872_inst_ack_1, ack => convTranspose_CP_772_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	159 
    -- CP-element group 160: 	127 
    -- CP-element group 160: 	131 
    -- CP-element group 160: 	135 
    -- CP-element group 160: 	139 
    -- CP-element group 160: 	143 
    -- CP-element group 160: 	147 
    -- CP-element group 160: 	151 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (9) 
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/word_access_start/word_0/rr
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/word_access_start/word_0/$entry
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/word_access_start/$entry
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/ptr_deref_880_Split/split_ack
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/ptr_deref_880_Split/split_req
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/ptr_deref_880_Split/$exit
      -- CP-element group 160: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/ptr_deref_880_Split/$entry
      -- 
    rr_2001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(160), ack => ptr_deref_880_store_0_req_0); -- 
    convTranspose_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(155) & convTranspose_CP_772_elements(159) & convTranspose_CP_772_elements(127) & convTranspose_CP_772_elements(131) & convTranspose_CP_772_elements(135) & convTranspose_CP_772_elements(139) & convTranspose_CP_772_elements(143) & convTranspose_CP_772_elements(147) & convTranspose_CP_772_elements(151);
      gj_convTranspose_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/word_access_start/word_0/ra
      -- CP-element group 161: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/word_access_start/word_0/$exit
      -- CP-element group 161: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/word_access_start/$exit
      -- CP-element group 161: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Sample/$exit
      -- 
    ra_2002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_880_store_0_ack_0, ack => convTranspose_CP_772_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	350 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/word_access_complete/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/word_access_complete/$exit
      -- CP-element group 162: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/word_access_complete/word_0/ca
      -- 
    ca_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_880_store_0_ack_1, ack => convTranspose_CP_772_elements(162)); -- 
    -- CP-element group 163:  branch  join  transition  place  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: 	124 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (10) 
      -- CP-element group 163: 	 branch_block_stmt_312/if_stmt_894_eval_test/$entry
      -- CP-element group 163: 	 branch_block_stmt_312/if_stmt_894_dead_link/$entry
      -- CP-element group 163: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893__exit__
      -- CP-element group 163: 	 branch_block_stmt_312/if_stmt_894__entry__
      -- CP-element group 163: 	 branch_block_stmt_312/if_stmt_894_eval_test/$exit
      -- CP-element group 163: 	 branch_block_stmt_312/R_exitcond32_895_place
      -- CP-element group 163: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/$exit
      -- CP-element group 163: 	 branch_block_stmt_312/if_stmt_894_else_link/$entry
      -- CP-element group 163: 	 branch_block_stmt_312/if_stmt_894_if_link/$entry
      -- CP-element group 163: 	 branch_block_stmt_312/if_stmt_894_eval_test/branch_req
      -- 
    branch_req_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(163), ack => if_stmt_894_branch_req_0); -- 
    convTranspose_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(162) & convTranspose_CP_772_elements(124);
      gj_convTranspose_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  merge  transition  place  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	344 
    -- CP-element group 164:  members (13) 
      -- CP-element group 164: 	 branch_block_stmt_312/merge_stmt_670__exit__
      -- CP-element group 164: 	 branch_block_stmt_312/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader
      -- CP-element group 164: 	 branch_block_stmt_312/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit
      -- CP-element group 164: 	 branch_block_stmt_312/if_stmt_894_if_link/if_choice_transition
      -- CP-element group 164: 	 branch_block_stmt_312/if_stmt_894_if_link/$exit
      -- CP-element group 164: 	 branch_block_stmt_312/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 164: 	 branch_block_stmt_312/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 164: 	 branch_block_stmt_312/merge_stmt_670_PhiReqMerge
      -- CP-element group 164: 	 branch_block_stmt_312/merge_stmt_670_PhiAck/$entry
      -- CP-element group 164: 	 branch_block_stmt_312/merge_stmt_670_PhiAck/$exit
      -- CP-element group 164: 	 branch_block_stmt_312/merge_stmt_670_PhiAck/dummy
      -- CP-element group 164: 	 branch_block_stmt_312/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader_PhiReq/$entry
      -- CP-element group 164: 	 branch_block_stmt_312/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_894_branch_ack_1, ack => convTranspose_CP_772_elements(164)); -- 
    -- CP-element group 165:  fork  transition  place  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	346 
    -- CP-element group 165: 	347 
    -- CP-element group 165:  members (12) 
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody
      -- CP-element group 165: 	 branch_block_stmt_312/if_stmt_894_else_link/else_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_312/if_stmt_894_else_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/$entry
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/$entry
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/$entry
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/$entry
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_894_branch_ack_0, ack => convTranspose_CP_772_elements(165)); -- 
    rr_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(165), ack => type_cast_735_inst_req_0); -- 
    cr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(165), ack => type_cast_735_inst_req_1); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	115 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_sample_completed_
      -- 
    ra_2044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_0, ack => convTranspose_CP_772_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	115 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	170 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_908_update_completed_
      -- 
    ca_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_1, ack => convTranspose_CP_772_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	115 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Sample/ra
      -- CP-element group 168: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_sample_completed_
      -- 
    ra_2058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_917_inst_ack_0, ack => convTranspose_CP_772_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	115 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/type_cast_917_update_completed_
      -- 
    ca_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_917_inst_ack_1, ack => convTranspose_CP_772_elements(169)); -- 
    -- CP-element group 170:  join  transition  place  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	167 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	351 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942__exit__
      -- CP-element group 170: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182
      -- CP-element group 170: 	 branch_block_stmt_312/assign_stmt_905_to_assign_stmt_942/$exit
      -- CP-element group 170: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/phi_stmt_945/$entry
      -- CP-element group 170: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/$entry
      -- 
    convTranspose_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(167) & convTranspose_CP_772_elements(169);
      gj_convTranspose_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	356 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	210 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Sample/ack
      -- CP-element group 171: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_sample_complete
      -- 
    ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_959_index_offset_ack_0, ack => convTranspose_CP_772_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	356 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (11) 
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_request/$entry
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_request/req
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_offset_calculated
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_sample_start_
      -- 
    ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_959_index_offset_ack_1, ack => convTranspose_CP_772_elements(172)); -- 
    req_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(172), ack => addr_of_960_final_reg_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_request/$exit
      -- CP-element group 173: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_request/ack
      -- CP-element group 173: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_sample_completed_
      -- 
    ack_2107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_960_final_reg_ack_0, ack => convTranspose_CP_772_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	356 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	207 
    -- CP-element group 174:  members (19) 
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_complete/ack
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_word_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_address_resized
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_addr_resize/$entry
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_addr_resize/$exit
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_addr_resize/base_resize_req
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_addr_resize/base_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_base_plus_offset/sum_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_word_addrgen/$entry
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_word_addrgen/$exit
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_word_addrgen/root_register_req
      -- CP-element group 174: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_word_addrgen/root_register_ack
      -- 
    ack_2112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_960_final_reg_ack_1, ack => convTranspose_CP_772_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	356 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_update_start_
      -- CP-element group 175: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_sample_completed_
      -- 
    ra_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_963_inst_ack_0, ack => convTranspose_CP_772_elements(175)); -- 
    cr_2125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(175), ack => RPIPE_ConvTranspose_input_pipe_963_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_update_completed_
      -- 
    ca_2126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_963_inst_ack_1, ack => convTranspose_CP_772_elements(176)); -- 
    rr_2134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(176), ack => type_cast_967_inst_req_0); -- 
    rr_2148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(176), ack => RPIPE_ConvTranspose_input_pipe_976_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_sample_completed_
      -- 
    ra_2135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_0, ack => convTranspose_CP_772_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	356 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	207 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_update_completed_
      -- 
    ca_2140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_1, ack => convTranspose_CP_772_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_update_start_
      -- CP-element group 179: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_sample_completed_
      -- 
    ra_2149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_976_inst_ack_0, ack => convTranspose_CP_772_elements(179)); -- 
    cr_2153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(179), ack => RPIPE_ConvTranspose_input_pipe_976_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_976_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_sample_start_
      -- 
    ca_2154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_976_inst_ack_1, ack => convTranspose_CP_772_elements(180)); -- 
    rr_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(180), ack => type_cast_980_inst_req_0); -- 
    rr_2176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(180), ack => RPIPE_ConvTranspose_input_pipe_994_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_sample_completed_
      -- 
    ra_2163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_980_inst_ack_0, ack => convTranspose_CP_772_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	356 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	207 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_update_completed_
      -- 
    ca_2168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_980_inst_ack_1, ack => convTranspose_CP_772_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_update_start_
      -- CP-element group 183: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_sample_completed_
      -- 
    ra_2177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_994_inst_ack_0, ack => convTranspose_CP_772_elements(183)); -- 
    cr_2181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(183), ack => RPIPE_ConvTranspose_input_pipe_994_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_994_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Sample/$entry
      -- 
    ca_2182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_994_inst_ack_1, ack => convTranspose_CP_772_elements(184)); -- 
    rr_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(184), ack => type_cast_998_inst_req_0); -- 
    rr_2204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(184), ack => RPIPE_ConvTranspose_input_pipe_1012_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_sample_completed_
      -- 
    ra_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_998_inst_ack_0, ack => convTranspose_CP_772_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	356 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	207 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Update/ca
      -- 
    ca_2196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_998_inst_ack_1, ack => convTranspose_CP_772_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_update_start_
      -- 
    ra_2205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1012_inst_ack_0, ack => convTranspose_CP_772_elements(187)); -- 
    cr_2209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(187), ack => RPIPE_ConvTranspose_input_pipe_1012_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1012_update_completed_
      -- 
    ca_2210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1012_inst_ack_1, ack => convTranspose_CP_772_elements(188)); -- 
    rr_2218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(188), ack => type_cast_1016_inst_req_0); -- 
    rr_2232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(188), ack => RPIPE_ConvTranspose_input_pipe_1030_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_sample_completed_
      -- 
    ra_2219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1016_inst_ack_0, ack => convTranspose_CP_772_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	356 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	207 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_update_completed_
      -- 
    ca_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1016_inst_ack_1, ack => convTranspose_CP_772_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_update_start_
      -- CP-element group 191: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_sample_completed_
      -- 
    ra_2233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1030_inst_ack_0, ack => convTranspose_CP_772_elements(191)); -- 
    cr_2237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(191), ack => RPIPE_ConvTranspose_input_pipe_1030_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1030_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_sample_start_
      -- 
    ca_2238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1030_inst_ack_1, ack => convTranspose_CP_772_elements(192)); -- 
    rr_2246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(192), ack => type_cast_1034_inst_req_0); -- 
    rr_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(192), ack => RPIPE_ConvTranspose_input_pipe_1048_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_sample_completed_
      -- 
    ra_2247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1034_inst_ack_0, ack => convTranspose_CP_772_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	356 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	207 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_update_completed_
      -- 
    ca_2252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1034_inst_ack_1, ack => convTranspose_CP_772_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_update_start_
      -- CP-element group 195: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Update/cr
      -- CP-element group 195: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Sample/ra
      -- 
    ra_2261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1048_inst_ack_0, ack => convTranspose_CP_772_elements(195)); -- 
    cr_2265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(195), ack => RPIPE_ConvTranspose_input_pipe_1048_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	199 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1048_Update/$exit
      -- 
    ca_2266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1048_inst_ack_1, ack => convTranspose_CP_772_elements(196)); -- 
    rr_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(196), ack => RPIPE_ConvTranspose_input_pipe_1066_inst_req_0); -- 
    rr_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(196), ack => type_cast_1052_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_sample_completed_
      -- 
    ra_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1052_inst_ack_0, ack => convTranspose_CP_772_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	356 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	207 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_update_completed_
      -- 
    ca_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1052_inst_ack_1, ack => convTranspose_CP_772_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_update_start_
      -- CP-element group 199: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Update/cr
      -- CP-element group 199: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Sample/$exit
      -- 
    ra_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1066_inst_ack_0, ack => convTranspose_CP_772_elements(199)); -- 
    cr_2293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(199), ack => RPIPE_ConvTranspose_input_pipe_1066_inst_req_1); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1066_update_completed_
      -- 
    ca_2294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1066_inst_ack_1, ack => convTranspose_CP_772_elements(200)); -- 
    rr_2302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(200), ack => type_cast_1070_inst_req_0); -- 
    rr_2316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(200), ack => RPIPE_ConvTranspose_input_pipe_1084_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Sample/ra
      -- 
    ra_2303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_0, ack => convTranspose_CP_772_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	356 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Update/$exit
      -- 
    ca_2308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_1, ack => convTranspose_CP_772_elements(202)); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Update/cr
      -- CP-element group 203: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_update_start_
      -- CP-element group 203: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Update/$entry
      -- 
    ra_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1084_inst_ack_0, ack => convTranspose_CP_772_elements(203)); -- 
    cr_2321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(203), ack => RPIPE_ConvTranspose_input_pipe_1084_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Sample/rr
      -- CP-element group 204: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_1084_Update/$exit
      -- 
    ca_2322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1084_inst_ack_1, ack => convTranspose_CP_772_elements(204)); -- 
    rr_2330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(204), ack => type_cast_1088_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Sample/ra
      -- CP-element group 205: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_sample_completed_
      -- 
    ra_2331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1088_inst_ack_0, ack => convTranspose_CP_772_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	356 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Update/ca
      -- 
    ca_2336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1088_inst_ack_1, ack => convTranspose_CP_772_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	198 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: 	174 
    -- CP-element group 207: 	178 
    -- CP-element group 207: 	182 
    -- CP-element group 207: 	186 
    -- CP-element group 207: 	190 
    -- CP-element group 207: 	194 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/ptr_deref_1096_Split/$entry
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/ptr_deref_1096_Split/$exit
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/ptr_deref_1096_Split/split_req
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/ptr_deref_1096_Split/split_ack
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/word_access_start/word_0/rr
      -- 
    rr_2374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(207), ack => ptr_deref_1096_store_0_req_0); -- 
    convTranspose_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(198) & convTranspose_CP_772_elements(202) & convTranspose_CP_772_elements(206) & convTranspose_CP_772_elements(174) & convTranspose_CP_772_elements(178) & convTranspose_CP_772_elements(182) & convTranspose_CP_772_elements(186) & convTranspose_CP_772_elements(190) & convTranspose_CP_772_elements(194);
      gj_convTranspose_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/word_access_start/$exit
      -- CP-element group 208: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/word_access_start/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Sample/word_access_start/word_0/ra
      -- 
    ra_2375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1096_store_0_ack_0, ack => convTranspose_CP_772_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	356 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/word_access_complete/$exit
      -- CP-element group 209: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/word_access_complete/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/word_access_complete/word_0/ca
      -- 
    ca_2386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1096_store_0_ack_1, ack => convTranspose_CP_772_elements(209)); -- 
    -- CP-element group 210:  branch  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: 	171 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (10) 
      -- CP-element group 210: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109__exit__
      -- CP-element group 210: 	 branch_block_stmt_312/if_stmt_1110__entry__
      -- CP-element group 210: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/$exit
      -- CP-element group 210: 	 branch_block_stmt_312/if_stmt_1110_dead_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_312/if_stmt_1110_eval_test/$entry
      -- CP-element group 210: 	 branch_block_stmt_312/if_stmt_1110_eval_test/$exit
      -- CP-element group 210: 	 branch_block_stmt_312/if_stmt_1110_eval_test/branch_req
      -- CP-element group 210: 	 branch_block_stmt_312/R_exitcond23_1111_place
      -- CP-element group 210: 	 branch_block_stmt_312/if_stmt_1110_if_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_312/if_stmt_1110_else_link/$entry
      -- 
    branch_req_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(210), ack => if_stmt_1110_branch_req_0); -- 
    convTranspose_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(209) & convTranspose_CP_772_elements(171);
      gj_convTranspose_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  transition  place  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	357 
    -- CP-element group 211:  members (13) 
      -- CP-element group 211: 	 branch_block_stmt_312/merge_stmt_1116__exit__
      -- CP-element group 211: 	 branch_block_stmt_312/forx_xend235x_xloopexit_forx_xend235
      -- CP-element group 211: 	 branch_block_stmt_312/if_stmt_1110_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_312/if_stmt_1110_if_link/if_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_312/forx_xbody182_forx_xend235x_xloopexit
      -- CP-element group 211: 	 branch_block_stmt_312/forx_xbody182_forx_xend235x_xloopexit_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_312/forx_xbody182_forx_xend235x_xloopexit_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_312/merge_stmt_1116_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_312/merge_stmt_1116_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_312/merge_stmt_1116_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_312/merge_stmt_1116_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_312/forx_xend235x_xloopexit_forx_xend235_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_312/forx_xend235x_xloopexit_forx_xend235_PhiReq/$exit
      -- 
    if_choice_transition_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1110_branch_ack_1, ack => convTranspose_CP_772_elements(211)); -- 
    -- CP-element group 212:  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	352 
    -- CP-element group 212: 	353 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_312/if_stmt_1110_else_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_312/if_stmt_1110_else_link/else_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/$entry
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/$entry
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/$entry
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1110_branch_ack_0, ack => convTranspose_CP_772_elements(212)); -- 
    rr_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(212), ack => type_cast_948_inst_req_0); -- 
    cr_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(212), ack => type_cast_948_inst_req_1); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	357 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Sample/ra
      -- 
    ra_2417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1121_inst_ack_0, ack => convTranspose_CP_772_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	357 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	219 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Update/ca
      -- 
    ca_2422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1121_inst_ack_1, ack => convTranspose_CP_772_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	357 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Sample/ra
      -- 
    ra_2431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1125_inst_ack_0, ack => convTranspose_CP_772_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	357 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	219 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Update/ca
      -- 
    ca_2436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1125_inst_ack_1, ack => convTranspose_CP_772_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	357 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Sample/ra
      -- 
    ra_2445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1129_inst_ack_0, ack => convTranspose_CP_772_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	357 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Update/ca
      -- 
    ca_2450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1129_inst_ack_1, ack => convTranspose_CP_772_elements(218)); -- 
    -- CP-element group 219:  branch  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	214 
    -- CP-element group 219: 	216 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (10) 
      -- CP-element group 219: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146__exit__
      -- CP-element group 219: 	 branch_block_stmt_312/if_stmt_1147__entry__
      -- CP-element group 219: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/$exit
      -- CP-element group 219: 	 branch_block_stmt_312/if_stmt_1147_dead_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_312/if_stmt_1147_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_312/if_stmt_1147_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_312/if_stmt_1147_eval_test/branch_req
      -- CP-element group 219: 	 branch_block_stmt_312/R_cmp249422_1148_place
      -- CP-element group 219: 	 branch_block_stmt_312/if_stmt_1147_if_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_312/if_stmt_1147_else_link/$entry
      -- 
    branch_req_2458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(219), ack => if_stmt_1147_branch_req_0); -- 
    convTranspose_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(214) & convTranspose_CP_772_elements(216) & convTranspose_CP_772_elements(218);
      gj_convTranspose_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: 	223 
    -- CP-element group 220: 	224 
    -- CP-element group 220: 	225 
    -- CP-element group 220: 	226 
    -- CP-element group 220: 	227 
    -- CP-element group 220:  members (30) 
      -- CP-element group 220: 	 branch_block_stmt_312/merge_stmt_1153__exit__
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194__entry__
      -- CP-element group 220: 	 branch_block_stmt_312/if_stmt_1147_if_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_312/if_stmt_1147_if_link/if_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_312/forx_xend235_bbx_xnph424
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_update_start_
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Update/cr
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_update_start_
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Update/cr
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_update_start_
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Update/cr
      -- CP-element group 220: 	 branch_block_stmt_312/forx_xend235_bbx_xnph424_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/forx_xend235_bbx_xnph424_PhiReq/$exit
      -- CP-element group 220: 	 branch_block_stmt_312/merge_stmt_1153_PhiReqMerge
      -- CP-element group 220: 	 branch_block_stmt_312/merge_stmt_1153_PhiAck/$entry
      -- CP-element group 220: 	 branch_block_stmt_312/merge_stmt_1153_PhiAck/$exit
      -- CP-element group 220: 	 branch_block_stmt_312/merge_stmt_1153_PhiAck/dummy
      -- 
    if_choice_transition_2463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1147_branch_ack_1, ack => convTranspose_CP_772_elements(220)); -- 
    rr_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(220), ack => type_cast_1156_inst_req_0); -- 
    cr_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(220), ack => type_cast_1156_inst_req_1); -- 
    rr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(220), ack => type_cast_1160_inst_req_0); -- 
    cr_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(220), ack => type_cast_1160_inst_req_1); -- 
    rr_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(220), ack => type_cast_1169_inst_req_0); -- 
    cr_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(220), ack => type_cast_1169_inst_req_1); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	364 
    -- CP-element group 221:  members (5) 
      -- CP-element group 221: 	 branch_block_stmt_312/if_stmt_1147_else_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_312/if_stmt_1147_else_link/else_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_312/forx_xend235_forx_xend257
      -- CP-element group 221: 	 branch_block_stmt_312/forx_xend235_forx_xend257_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_312/forx_xend235_forx_xend257_PhiReq/$exit
      -- 
    else_choice_transition_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1147_branch_ack_0, ack => convTranspose_CP_772_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_sample_completed_
      -- CP-element group 222: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Sample/ra
      -- 
    ra_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_0, ack => convTranspose_CP_772_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	228 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1156_Update/ca
      -- 
    ca_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_1, ack => convTranspose_CP_772_elements(223)); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	220 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Sample/ra
      -- 
    ra_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_0, ack => convTranspose_CP_772_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	220 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	228 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1160_Update/ca
      -- 
    ca_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_1, ack => convTranspose_CP_772_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	220 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Sample/ra
      -- 
    ra_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_0, ack => convTranspose_CP_772_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	220 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/type_cast_1169_Update/ca
      -- 
    ca_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_1, ack => convTranspose_CP_772_elements(227)); -- 
    -- CP-element group 228:  join  transition  place  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	223 
    -- CP-element group 228: 	225 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	358 
    -- CP-element group 228:  members (6) 
      -- CP-element group 228: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194__exit__
      -- CP-element group 228: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251
      -- CP-element group 228: 	 branch_block_stmt_312/assign_stmt_1157_to_assign_stmt_1194/$exit
      -- CP-element group 228: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/phi_stmt_1197/$entry
      -- CP-element group 228: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/$entry
      -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(223) & convTranspose_CP_772_elements(225) & convTranspose_CP_772_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	363 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	235 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_sample_complete
      -- CP-element group 229: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Sample/ack
      -- 
    ack_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1211_index_offset_ack_0, ack => convTranspose_CP_772_elements(229)); -- 
    -- CP-element group 230:  transition  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	363 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (11) 
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_root_address_calculated
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_offset_calculated
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Update/ack
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_base_plus_offset/$entry
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_base_plus_offset/$exit
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_base_plus_offset/sum_rename_req
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_base_plus_offset/sum_rename_ack
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_request/$entry
      -- CP-element group 230: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_request/req
      -- 
    ack_2548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1211_index_offset_ack_1, ack => convTranspose_CP_772_elements(230)); -- 
    req_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(230), ack => addr_of_1212_final_reg_req_0); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_request/$exit
      -- CP-element group 231: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_request/ack
      -- 
    ack_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1212_final_reg_ack_0, ack => convTranspose_CP_772_elements(231)); -- 
    -- CP-element group 232:  join  fork  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	363 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (28) 
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_complete/$exit
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_complete/ack
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_word_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_root_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_address_resized
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_addr_resize/$entry
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_addr_resize/$exit
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_addr_resize/base_resize_req
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_addr_resize/base_resize_ack
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_plus_offset/$entry
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_plus_offset/$exit
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_plus_offset/sum_rename_req
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_base_plus_offset/sum_rename_ack
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_word_addrgen/$entry
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_word_addrgen/$exit
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_word_addrgen/root_register_req
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_word_addrgen/root_register_ack
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/ptr_deref_1215_Split/$entry
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/ptr_deref_1215_Split/$exit
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/ptr_deref_1215_Split/split_req
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/ptr_deref_1215_Split/split_ack
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/word_access_start/$entry
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/word_access_start/word_0/$entry
      -- CP-element group 232: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/word_access_start/word_0/rr
      -- 
    ack_2563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1212_final_reg_ack_1, ack => convTranspose_CP_772_elements(232)); -- 
    rr_2601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(232), ack => ptr_deref_1215_store_0_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (5) 
      -- CP-element group 233: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/word_access_start/$exit
      -- CP-element group 233: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/word_access_start/word_0/$exit
      -- CP-element group 233: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Sample/word_access_start/word_0/ra
      -- 
    ra_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1215_store_0_ack_0, ack => convTranspose_CP_772_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	363 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (5) 
      -- CP-element group 234: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/word_access_complete/$exit
      -- CP-element group 234: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/word_access_complete/word_0/$exit
      -- CP-element group 234: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/word_access_complete/word_0/ca
      -- 
    ca_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1215_store_0_ack_1, ack => convTranspose_CP_772_elements(234)); -- 
    -- CP-element group 235:  branch  join  transition  place  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	229 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (10) 
      -- CP-element group 235: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229__exit__
      -- CP-element group 235: 	 branch_block_stmt_312/if_stmt_1230__entry__
      -- CP-element group 235: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/$exit
      -- CP-element group 235: 	 branch_block_stmt_312/if_stmt_1230_dead_link/$entry
      -- CP-element group 235: 	 branch_block_stmt_312/if_stmt_1230_eval_test/$entry
      -- CP-element group 235: 	 branch_block_stmt_312/if_stmt_1230_eval_test/$exit
      -- CP-element group 235: 	 branch_block_stmt_312/if_stmt_1230_eval_test/branch_req
      -- CP-element group 235: 	 branch_block_stmt_312/R_exitcond_1231_place
      -- CP-element group 235: 	 branch_block_stmt_312/if_stmt_1230_if_link/$entry
      -- CP-element group 235: 	 branch_block_stmt_312/if_stmt_1230_else_link/$entry
      -- 
    branch_req_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(235), ack => if_stmt_1230_branch_req_0); -- 
    convTranspose_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(229) & convTranspose_CP_772_elements(234);
      gj_convTranspose_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  merge  transition  place  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	364 
    -- CP-element group 236:  members (13) 
      -- CP-element group 236: 	 branch_block_stmt_312/merge_stmt_1236__exit__
      -- CP-element group 236: 	 branch_block_stmt_312/forx_xend257x_xloopexit_forx_xend257
      -- CP-element group 236: 	 branch_block_stmt_312/if_stmt_1230_if_link/$exit
      -- CP-element group 236: 	 branch_block_stmt_312/if_stmt_1230_if_link/if_choice_transition
      -- CP-element group 236: 	 branch_block_stmt_312/forx_xbody251_forx_xend257x_xloopexit
      -- CP-element group 236: 	 branch_block_stmt_312/forx_xbody251_forx_xend257x_xloopexit_PhiReq/$entry
      -- CP-element group 236: 	 branch_block_stmt_312/forx_xbody251_forx_xend257x_xloopexit_PhiReq/$exit
      -- CP-element group 236: 	 branch_block_stmt_312/merge_stmt_1236_PhiReqMerge
      -- CP-element group 236: 	 branch_block_stmt_312/merge_stmt_1236_PhiAck/$entry
      -- CP-element group 236: 	 branch_block_stmt_312/merge_stmt_1236_PhiAck/$exit
      -- CP-element group 236: 	 branch_block_stmt_312/merge_stmt_1236_PhiAck/dummy
      -- CP-element group 236: 	 branch_block_stmt_312/forx_xend257x_xloopexit_forx_xend257_PhiReq/$entry
      -- CP-element group 236: 	 branch_block_stmt_312/forx_xend257x_xloopexit_forx_xend257_PhiReq/$exit
      -- 
    if_choice_transition_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1230_branch_ack_1, ack => convTranspose_CP_772_elements(236)); -- 
    -- CP-element group 237:  fork  transition  place  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	359 
    -- CP-element group 237: 	360 
    -- CP-element group 237:  members (12) 
      -- CP-element group 237: 	 branch_block_stmt_312/if_stmt_1230_else_link/$exit
      -- CP-element group 237: 	 branch_block_stmt_312/if_stmt_1230_else_link/else_choice_transition
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/$entry
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/$entry
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/$entry
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/$entry
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/$entry
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Sample/rr
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1230_branch_ack_0, ack => convTranspose_CP_772_elements(237)); -- 
    rr_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(237), ack => type_cast_1203_inst_req_0); -- 
    cr_3545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(237), ack => type_cast_1203_inst_req_1); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	364 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Sample/cra
      -- 
    cra_2644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1241_call_ack_0, ack => convTranspose_CP_772_elements(238)); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	364 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Update/cca
      -- CP-element group 239: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Sample/rr
      -- 
    cca_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1241_call_ack_1, ack => convTranspose_CP_772_elements(239)); -- 
    rr_2657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(239), ack => type_cast_1246_inst_req_0); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Sample/ra
      -- 
    ra_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_0, ack => convTranspose_CP_772_elements(240)); -- 
    -- CP-element group 241:  fork  transition  place  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	364 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (13) 
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247__exit__
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263__entry__
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/$exit
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Update/ca
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263/$entry
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_update_start_
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Sample/crr
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Update/ccr
      -- 
    ca_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_1, ack => convTranspose_CP_772_elements(241)); -- 
    crr_2674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(241), ack => call_stmt_1263_call_req_0); -- 
    ccr_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(241), ack => call_stmt_1263_call_req_1); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Sample/cra
      -- 
    cra_2675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1263_call_ack_0, ack => convTranspose_CP_772_elements(242)); -- 
    -- CP-element group 243:  fork  transition  place  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: 	245 
    -- CP-element group 243: 	247 
    -- CP-element group 243:  members (16) 
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1263__exit__
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276__entry__
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1263/$exit
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1263/call_stmt_1263_Update/cca
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/$entry
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_update_start_
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Sample/crr
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Update/ccr
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_update_start_
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Update/cr
      -- 
    cca_2680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1263_call_ack_1, ack => convTranspose_CP_772_elements(243)); -- 
    crr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(243), ack => call_stmt_1266_call_req_0); -- 
    ccr_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(243), ack => call_stmt_1266_call_req_1); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(243), ack => type_cast_1270_inst_req_1); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Sample/cra
      -- 
    cra_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1266_call_ack_0, ack => convTranspose_CP_772_elements(244)); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/call_stmt_1266_Update/cca
      -- CP-element group 245: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Sample/rr
      -- 
    cca_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1266_call_ack_1, ack => convTranspose_CP_772_elements(245)); -- 
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(245), ack => type_cast_1270_inst_req_0); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Sample/ra
      -- 
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_0, ack => convTranspose_CP_772_elements(246)); -- 
    -- CP-element group 247:  fork  transition  place  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	243 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247: 	249 
    -- CP-element group 247: 	250 
    -- CP-element group 247: 	251 
    -- CP-element group 247: 	252 
    -- CP-element group 247: 	253 
    -- CP-element group 247: 	254 
    -- CP-element group 247: 	255 
    -- CP-element group 247: 	256 
    -- CP-element group 247: 	257 
    -- CP-element group 247: 	258 
    -- CP-element group 247: 	259 
    -- CP-element group 247: 	260 
    -- CP-element group 247: 	261 
    -- CP-element group 247: 	262 
    -- CP-element group 247: 	263 
    -- CP-element group 247:  members (55) 
      -- CP-element group 247: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276__exit__
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375__entry__
      -- CP-element group 247: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/$exit
      -- CP-element group 247: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_312/call_stmt_1266_to_assign_stmt_1276/type_cast_1270_Update/ca
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_update_start_
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Update/cr
      -- 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_1, ack => convTranspose_CP_772_elements(247)); -- 
    rr_2722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1280_inst_req_0); -- 
    cr_2727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1280_inst_req_1); -- 
    rr_2736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1290_inst_req_0); -- 
    cr_2741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1290_inst_req_1); -- 
    rr_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1300_inst_req_0); -- 
    cr_2755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1300_inst_req_1); -- 
    rr_2764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1310_inst_req_0); -- 
    cr_2769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1310_inst_req_1); -- 
    rr_2778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1320_inst_req_0); -- 
    cr_2783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1320_inst_req_1); -- 
    rr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1330_inst_req_0); -- 
    cr_2797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1330_inst_req_1); -- 
    rr_2806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1340_inst_req_0); -- 
    cr_2811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1340_inst_req_1); -- 
    rr_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1350_inst_req_0); -- 
    cr_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(247), ack => type_cast_1350_inst_req_1); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Sample/ra
      -- 
    ra_2723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1280_inst_ack_0, ack => convTranspose_CP_772_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	284 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1280_Update/ca
      -- 
    ca_2728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1280_inst_ack_1, ack => convTranspose_CP_772_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	247 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Sample/ra
      -- 
    ra_2737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1290_inst_ack_0, ack => convTranspose_CP_772_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	247 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	281 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1290_Update/ca
      -- 
    ca_2742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1290_inst_ack_1, ack => convTranspose_CP_772_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	247 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Sample/ra
      -- 
    ra_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_0, ack => convTranspose_CP_772_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	247 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	278 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1300_Update/ca
      -- 
    ca_2756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_1, ack => convTranspose_CP_772_elements(253)); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	247 
    -- CP-element group 254: successors 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Sample/ra
      -- 
    ra_2765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_0, ack => convTranspose_CP_772_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	247 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	275 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1310_Update/ca
      -- 
    ca_2770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_1, ack => convTranspose_CP_772_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	247 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Sample/ra
      -- 
    ra_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_0, ack => convTranspose_CP_772_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	247 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	272 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1320_Update/ca
      -- 
    ca_2784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_1, ack => convTranspose_CP_772_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	247 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Sample/ra
      -- 
    ra_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1330_inst_ack_0, ack => convTranspose_CP_772_elements(258)); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	247 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	269 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1330_Update/ca
      -- 
    ca_2798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1330_inst_ack_1, ack => convTranspose_CP_772_elements(259)); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	247 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Sample/ra
      -- 
    ra_2807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1340_inst_ack_0, ack => convTranspose_CP_772_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	247 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	266 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1340_Update/ca
      -- 
    ca_2812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1340_inst_ack_1, ack => convTranspose_CP_772_elements(261)); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	247 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Sample/ra
      -- 
    ra_2821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1350_inst_ack_0, ack => convTranspose_CP_772_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	247 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/type_cast_1350_Update/ca
      -- CP-element group 263: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Sample/req
      -- 
    ca_2826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1350_inst_ack_1, ack => convTranspose_CP_772_elements(263)); -- 
    req_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(263), ack => WPIPE_ConvTranspose_output_pipe_1352_inst_req_0); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_update_start_
      -- CP-element group 264: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Sample/ack
      -- CP-element group 264: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Update/req
      -- 
    ack_2835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1352_inst_ack_0, ack => convTranspose_CP_772_elements(264)); -- 
    req_2839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(264), ack => WPIPE_ConvTranspose_output_pipe_1352_inst_req_1); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1352_Update/ack
      -- 
    ack_2840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1352_inst_ack_1, ack => convTranspose_CP_772_elements(265)); -- 
    -- CP-element group 266:  join  transition  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	261 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Sample/req
      -- 
    req_2848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(266), ack => WPIPE_ConvTranspose_output_pipe_1355_inst_req_0); -- 
    convTranspose_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(261) & convTranspose_CP_772_elements(265);
      gj_convTranspose_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Update/req
      -- CP-element group 267: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_update_start_
      -- CP-element group 267: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Sample/ack
      -- 
    ack_2849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1355_inst_ack_0, ack => convTranspose_CP_772_elements(267)); -- 
    req_2853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(267), ack => WPIPE_ConvTranspose_output_pipe_1355_inst_req_1); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1355_update_completed_
      -- 
    ack_2854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1355_inst_ack_1, ack => convTranspose_CP_772_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	259 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Sample/req
      -- 
    req_2862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(269), ack => WPIPE_ConvTranspose_output_pipe_1358_inst_req_0); -- 
    convTranspose_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(259) & convTranspose_CP_772_elements(268);
      gj_convTranspose_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_update_start_
      -- CP-element group 270: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Update/req
      -- CP-element group 270: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Sample/ack
      -- 
    ack_2863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1358_inst_ack_0, ack => convTranspose_CP_772_elements(270)); -- 
    req_2867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(270), ack => WPIPE_ConvTranspose_output_pipe_1358_inst_req_1); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Update/ack
      -- CP-element group 271: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1358_Update/$exit
      -- 
    ack_2868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1358_inst_ack_1, ack => convTranspose_CP_772_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	257 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_sample_start_
      -- 
    req_2876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(272), ack => WPIPE_ConvTranspose_output_pipe_1361_inst_req_0); -- 
    convTranspose_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(257) & convTranspose_CP_772_elements(271);
      gj_convTranspose_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Update/req
      -- CP-element group 273: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_update_start_
      -- CP-element group 273: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_sample_completed_
      -- 
    ack_2877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1361_inst_ack_0, ack => convTranspose_CP_772_elements(273)); -- 
    req_2881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(273), ack => WPIPE_ConvTranspose_output_pipe_1361_inst_req_1); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1361_Update/ack
      -- 
    ack_2882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1361_inst_ack_1, ack => convTranspose_CP_772_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	255 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Sample/req
      -- CP-element group 275: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_sample_start_
      -- 
    req_2890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(275), ack => WPIPE_ConvTranspose_output_pipe_1364_inst_req_0); -- 
    convTranspose_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(255) & convTranspose_CP_772_elements(274);
      gj_convTranspose_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_update_start_
      -- CP-element group 276: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Sample/ack
      -- CP-element group 276: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Update/req
      -- CP-element group 276: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Update/$entry
      -- 
    ack_2891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1364_inst_ack_0, ack => convTranspose_CP_772_elements(276)); -- 
    req_2895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(276), ack => WPIPE_ConvTranspose_output_pipe_1364_inst_req_1); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Update/ack
      -- CP-element group 277: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1364_Update/$exit
      -- 
    ack_2896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1364_inst_ack_1, ack => convTranspose_CP_772_elements(277)); -- 
    -- CP-element group 278:  join  transition  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	253 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_sample_start_
      -- 
    req_2904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(278), ack => WPIPE_ConvTranspose_output_pipe_1367_inst_req_0); -- 
    convTranspose_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(253) & convTranspose_CP_772_elements(277);
      gj_convTranspose_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_update_start_
      -- CP-element group 279: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Update/req
      -- CP-element group 279: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Update/$entry
      -- 
    ack_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1367_inst_ack_0, ack => convTranspose_CP_772_elements(279)); -- 
    req_2909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(279), ack => WPIPE_ConvTranspose_output_pipe_1367_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1367_Update/$exit
      -- 
    ack_2910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1367_inst_ack_1, ack => convTranspose_CP_772_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	251 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Sample/req
      -- CP-element group 281: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_sample_start_
      -- 
    req_2918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(281), ack => WPIPE_ConvTranspose_output_pipe_1370_inst_req_0); -- 
    convTranspose_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(251) & convTranspose_CP_772_elements(280);
      gj_convTranspose_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Update/req
      -- CP-element group 282: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Update/$entry
      -- CP-element group 282: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Sample/ack
      -- CP-element group 282: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_update_start_
      -- CP-element group 282: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_sample_completed_
      -- 
    ack_2919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1370_inst_ack_0, ack => convTranspose_CP_772_elements(282)); -- 
    req_2923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(282), ack => WPIPE_ConvTranspose_output_pipe_1370_inst_req_1); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Update/ack
      -- CP-element group 283: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1370_update_completed_
      -- 
    ack_2924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1370_inst_ack_1, ack => convTranspose_CP_772_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	249 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Sample/req
      -- CP-element group 284: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_sample_start_
      -- 
    req_2932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(284), ack => WPIPE_ConvTranspose_output_pipe_1373_inst_req_0); -- 
    convTranspose_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(249) & convTranspose_CP_772_elements(283);
      gj_convTranspose_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Update/req
      -- CP-element group 285: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_update_start_
      -- CP-element group 285: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_sample_completed_
      -- 
    ack_2933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1373_inst_ack_0, ack => convTranspose_CP_772_elements(285)); -- 
    req_2937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(285), ack => WPIPE_ConvTranspose_output_pipe_1373_inst_req_1); -- 
    -- CP-element group 286:  branch  transition  place  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (13) 
      -- CP-element group 286: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375__exit__
      -- CP-element group 286: 	 branch_block_stmt_312/if_stmt_1377__entry__
      -- CP-element group 286: 	 branch_block_stmt_312/if_stmt_1377_else_link/$entry
      -- CP-element group 286: 	 branch_block_stmt_312/if_stmt_1377_if_link/$entry
      -- CP-element group 286: 	 branch_block_stmt_312/if_stmt_1377_eval_test/branch_req
      -- CP-element group 286: 	 branch_block_stmt_312/if_stmt_1377_eval_test/$exit
      -- CP-element group 286: 	 branch_block_stmt_312/if_stmt_1377_eval_test/$entry
      -- CP-element group 286: 	 branch_block_stmt_312/if_stmt_1377_dead_link/$entry
      -- CP-element group 286: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/WPIPE_ConvTranspose_output_pipe_1373_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_312/assign_stmt_1281_to_assign_stmt_1375/$exit
      -- CP-element group 286: 	 branch_block_stmt_312/R_cmp249422_1378_place
      -- 
    ack_2938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1373_inst_ack_1, ack => convTranspose_CP_772_elements(286)); -- 
    branch_req_2946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(286), ack => if_stmt_1377_branch_req_0); -- 
    -- CP-element group 287:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	289 
    -- CP-element group 287: 	290 
    -- CP-element group 287: 	291 
    -- CP-element group 287: 	292 
    -- CP-element group 287: 	293 
    -- CP-element group 287: 	294 
    -- CP-element group 287:  members (30) 
      -- CP-element group 287: 	 branch_block_stmt_312/merge_stmt_1383__exit__
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424__entry__
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_update_start_
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/if_stmt_1377_if_link/if_choice_transition
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_312/if_stmt_1377_if_link/$exit
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_update_start_
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_update_start_
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_312/forx_xend257_bbx_xnph
      -- CP-element group 287: 	 branch_block_stmt_312/forx_xend257_bbx_xnph_PhiReq/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/forx_xend257_bbx_xnph_PhiReq/$exit
      -- CP-element group 287: 	 branch_block_stmt_312/merge_stmt_1383_PhiReqMerge
      -- CP-element group 287: 	 branch_block_stmt_312/merge_stmt_1383_PhiAck/$entry
      -- CP-element group 287: 	 branch_block_stmt_312/merge_stmt_1383_PhiAck/$exit
      -- CP-element group 287: 	 branch_block_stmt_312/merge_stmt_1383_PhiAck/dummy
      -- 
    if_choice_transition_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1377_branch_ack_1, ack => convTranspose_CP_772_elements(287)); -- 
    rr_2968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(287), ack => type_cast_1386_inst_req_0); -- 
    cr_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(287), ack => type_cast_1399_inst_req_1); -- 
    rr_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(287), ack => type_cast_1399_inst_req_0); -- 
    cr_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(287), ack => type_cast_1390_inst_req_1); -- 
    rr_2982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(287), ack => type_cast_1390_inst_req_0); -- 
    cr_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(287), ack => type_cast_1386_inst_req_1); -- 
    -- CP-element group 288:  transition  place  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	371 
    -- CP-element group 288:  members (5) 
      -- CP-element group 288: 	 branch_block_stmt_312/if_stmt_1377_else_link/else_choice_transition
      -- CP-element group 288: 	 branch_block_stmt_312/if_stmt_1377_else_link/$exit
      -- CP-element group 288: 	 branch_block_stmt_312/forx_xend257_forx_xend417
      -- CP-element group 288: 	 branch_block_stmt_312/forx_xend257_forx_xend417_PhiReq/$entry
      -- CP-element group 288: 	 branch_block_stmt_312/forx_xend257_forx_xend417_PhiReq/$exit
      -- 
    else_choice_transition_2955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1377_branch_ack_0, ack => convTranspose_CP_772_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_sample_completed_
      -- CP-element group 289: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Sample/ra
      -- 
    ra_2969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_0, ack => convTranspose_CP_772_elements(289)); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	287 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	295 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Update/ca
      -- CP-element group 290: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1386_Update/$exit
      -- 
    ca_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_1, ack => convTranspose_CP_772_elements(290)); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	287 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Sample/ra
      -- CP-element group 291: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_sample_completed_
      -- 
    ra_2983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1390_inst_ack_0, ack => convTranspose_CP_772_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	287 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	295 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Update/ca
      -- CP-element group 292: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1390_update_completed_
      -- 
    ca_2988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1390_inst_ack_1, ack => convTranspose_CP_772_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	287 
    -- CP-element group 293: successors 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Sample/ra
      -- CP-element group 293: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_sample_completed_
      -- 
    ra_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_0, ack => convTranspose_CP_772_elements(293)); -- 
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	287 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Update/ca
      -- CP-element group 294: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/type_cast_1399_update_completed_
      -- 
    ca_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_1, ack => convTranspose_CP_772_elements(294)); -- 
    -- CP-element group 295:  join  transition  place  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	290 
    -- CP-element group 295: 	292 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	365 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424/$exit
      -- CP-element group 295: 	 branch_block_stmt_312/assign_stmt_1387_to_assign_stmt_1424__exit__
      -- CP-element group 295: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345
      -- CP-element group 295: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/$entry
      -- CP-element group 295: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/phi_stmt_1427/$entry
      -- CP-element group 295: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$entry
      -- 
    convTranspose_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(290) & convTranspose_CP_772_elements(292) & convTranspose_CP_772_elements(294);
      gj_convTranspose_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	370 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	341 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Sample/ack
      -- CP-element group 296: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_sample_complete
      -- 
    ack_3031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_index_offset_ack_0, ack => convTranspose_CP_772_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	370 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (11) 
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_root_address_calculated
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_offset_calculated
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_request/req
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_request/$entry
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_base_plus_offset/sum_rename_ack
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_base_plus_offset/sum_rename_req
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_base_plus_offset/$exit
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_base_plus_offset/$entry
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Update/ack
      -- CP-element group 297: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Update/$exit
      -- 
    ack_3036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_index_offset_ack_1, ack => convTranspose_CP_772_elements(297)); -- 
    req_3045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(297), ack => addr_of_1442_final_reg_req_0); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_sample_completed_
      -- CP-element group 298: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_request/ack
      -- CP-element group 298: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_request/$exit
      -- 
    ack_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1442_final_reg_ack_0, ack => convTranspose_CP_772_elements(298)); -- 
    -- CP-element group 299:  join  fork  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	370 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (24) 
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_update_completed_
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_word_addrgen/root_register_ack
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_word_addrgen/root_register_req
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_word_addrgen/$exit
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_word_addrgen/$entry
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_plus_offset/sum_rename_ack
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_plus_offset/sum_rename_req
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_plus_offset/$exit
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_plus_offset/$entry
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_addr_resize/base_resize_ack
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_addr_resize/base_resize_req
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_addr_resize/$exit
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_addr_resize/$entry
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_address_resized
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_root_address_calculated
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_word_address_calculated
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_base_address_calculated
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_sample_start_
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_complete/ack
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_complete/$exit
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/word_access_start/word_0/rr
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/word_access_start/word_0/$entry
      -- CP-element group 299: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/word_access_start/$entry
      -- 
    ack_3051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1442_final_reg_ack_1, ack => convTranspose_CP_772_elements(299)); -- 
    rr_3084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(299), ack => ptr_deref_1446_load_0_req_0); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300:  members (5) 
      -- CP-element group 300: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/word_access_start/word_0/ra
      -- CP-element group 300: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/word_access_start/word_0/$exit
      -- CP-element group 300: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Sample/word_access_start/$exit
      -- 
    ra_3085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1446_load_0_ack_0, ack => convTranspose_CP_772_elements(300)); -- 
    -- CP-element group 301:  fork  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	370 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301: 	304 
    -- CP-element group 301: 	306 
    -- CP-element group 301: 	308 
    -- CP-element group 301: 	310 
    -- CP-element group 301: 	312 
    -- CP-element group 301: 	314 
    -- CP-element group 301: 	316 
    -- CP-element group 301:  members (33) 
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/ptr_deref_1446_Merge/merge_ack
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/ptr_deref_1446_Merge/merge_req
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/ptr_deref_1446_Merge/$exit
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/ptr_deref_1446_Merge/$entry
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/word_access_complete/word_0/ca
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/word_access_complete/word_0/$exit
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/word_access_complete/$exit
      -- CP-element group 301: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/$exit
      -- 
    ca_3096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1446_load_0_ack_1, ack => convTranspose_CP_772_elements(301)); -- 
    rr_3109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1450_inst_req_0); -- 
    rr_3123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1460_inst_req_0); -- 
    rr_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1470_inst_req_0); -- 
    rr_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1480_inst_req_0); -- 
    rr_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1490_inst_req_0); -- 
    rr_3179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1500_inst_req_0); -- 
    rr_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1510_inst_req_0); -- 
    rr_3207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(301), ack => type_cast_1520_inst_req_0); -- 
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Sample/ra
      -- CP-element group 302: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Sample/$exit
      -- CP-element group 302: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_sample_completed_
      -- 
    ra_3110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1450_inst_ack_0, ack => convTranspose_CP_772_elements(302)); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	370 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	338 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Update/ca
      -- CP-element group 303: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Update/$exit
      -- CP-element group 303: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_update_completed_
      -- 
    ca_3115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1450_inst_ack_1, ack => convTranspose_CP_772_elements(303)); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	301 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Sample/ra
      -- CP-element group 304: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_sample_completed_
      -- 
    ra_3124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1460_inst_ack_0, ack => convTranspose_CP_772_elements(304)); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	370 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	335 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Update/ca
      -- CP-element group 305: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Update/$exit
      -- CP-element group 305: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_update_completed_
      -- 
    ca_3129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1460_inst_ack_1, ack => convTranspose_CP_772_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	301 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Sample/ra
      -- CP-element group 306: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_sample_completed_
      -- 
    ra_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1470_inst_ack_0, ack => convTranspose_CP_772_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	370 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	332 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Update/ca
      -- CP-element group 307: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_update_completed_
      -- 
    ca_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1470_inst_ack_1, ack => convTranspose_CP_772_elements(307)); -- 
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	301 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Sample/ra
      -- CP-element group 308: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Sample/$exit
      -- CP-element group 308: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_sample_completed_
      -- 
    ra_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1480_inst_ack_0, ack => convTranspose_CP_772_elements(308)); -- 
    -- CP-element group 309:  transition  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	370 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	329 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Update/ca
      -- CP-element group 309: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_update_completed_
      -- 
    ca_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1480_inst_ack_1, ack => convTranspose_CP_772_elements(309)); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	301 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Sample/ra
      -- CP-element group 310: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Sample/$exit
      -- 
    ra_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1490_inst_ack_0, ack => convTranspose_CP_772_elements(310)); -- 
    -- CP-element group 311:  transition  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	370 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	326 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Update/ca
      -- CP-element group 311: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Update/$exit
      -- 
    ca_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1490_inst_ack_1, ack => convTranspose_CP_772_elements(311)); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	301 
    -- CP-element group 312: successors 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Sample/ra
      -- 
    ra_3180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1500_inst_ack_0, ack => convTranspose_CP_772_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	370 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	323 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Update/ca
      -- CP-element group 313: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Update/$exit
      -- 
    ca_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1500_inst_ack_1, ack => convTranspose_CP_772_elements(313)); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	301 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Sample/ra
      -- CP-element group 314: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_sample_completed_
      -- 
    ra_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_0, ack => convTranspose_CP_772_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	370 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	320 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Update/ca
      -- CP-element group 315: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Update/$exit
      -- CP-element group 315: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_update_completed_
      -- 
    ca_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_1, ack => convTranspose_CP_772_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	301 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_sample_completed_
      -- CP-element group 316: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Sample/ra
      -- 
    ra_3208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1520_inst_ack_0, ack => convTranspose_CP_772_elements(316)); -- 
    -- CP-element group 317:  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	370 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_update_completed_
      -- CP-element group 317: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Sample/req
      -- CP-element group 317: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Update/ca
      -- CP-element group 317: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Update/$exit
      -- 
    ca_3213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1520_inst_ack_1, ack => convTranspose_CP_772_elements(317)); -- 
    req_3221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(317), ack => WPIPE_ConvTranspose_output_pipe_1522_inst_req_0); -- 
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Update/req
      -- CP-element group 318: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_update_start_
      -- CP-element group 318: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_sample_completed_
      -- 
    ack_3222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1522_inst_ack_0, ack => convTranspose_CP_772_elements(318)); -- 
    req_3226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(318), ack => WPIPE_ConvTranspose_output_pipe_1522_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Update/ack
      -- CP-element group 319: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1522_update_completed_
      -- 
    ack_3227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1522_inst_ack_1, ack => convTranspose_CP_772_elements(319)); -- 
    -- CP-element group 320:  join  transition  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	315 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Sample/req
      -- CP-element group 320: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_sample_start_
      -- 
    req_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(320), ack => WPIPE_ConvTranspose_output_pipe_1525_inst_req_0); -- 
    convTranspose_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(315) & convTranspose_CP_772_elements(319);
      gj_convTranspose_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Update/req
      -- CP-element group 321: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Sample/ack
      -- CP-element group 321: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_update_start_
      -- CP-element group 321: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_sample_completed_
      -- 
    ack_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1525_inst_ack_0, ack => convTranspose_CP_772_elements(321)); -- 
    req_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(321), ack => WPIPE_ConvTranspose_output_pipe_1525_inst_req_1); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Update/ack
      -- CP-element group 322: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1525_update_completed_
      -- 
    ack_3241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1525_inst_ack_1, ack => convTranspose_CP_772_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	313 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Sample/req
      -- CP-element group 323: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_sample_start_
      -- 
    req_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(323), ack => WPIPE_ConvTranspose_output_pipe_1528_inst_req_0); -- 
    convTranspose_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(313) & convTranspose_CP_772_elements(322);
      gj_convTranspose_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Sample/ack
      -- CP-element group 324: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Update/$entry
      -- CP-element group 324: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Update/req
      -- CP-element group 324: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_update_start_
      -- CP-element group 324: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_sample_completed_
      -- 
    ack_3250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1528_inst_ack_0, ack => convTranspose_CP_772_elements(324)); -- 
    req_3254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(324), ack => WPIPE_ConvTranspose_output_pipe_1528_inst_req_1); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1528_Update/ack
      -- 
    ack_3255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1528_inst_ack_1, ack => convTranspose_CP_772_elements(325)); -- 
    -- CP-element group 326:  join  transition  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	311 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Sample/req
      -- CP-element group 326: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_sample_start_
      -- 
    req_3263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(326), ack => WPIPE_ConvTranspose_output_pipe_1531_inst_req_0); -- 
    convTranspose_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(311) & convTranspose_CP_772_elements(325);
      gj_convTranspose_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_update_start_
      -- CP-element group 327: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Update/req
      -- CP-element group 327: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Update/$entry
      -- 
    ack_3264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1531_inst_ack_0, ack => convTranspose_CP_772_elements(327)); -- 
    req_3268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(327), ack => WPIPE_ConvTranspose_output_pipe_1531_inst_req_1); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1531_Update/$exit
      -- 
    ack_3269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1531_inst_ack_1, ack => convTranspose_CP_772_elements(328)); -- 
    -- CP-element group 329:  join  transition  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	309 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Sample/req
      -- CP-element group 329: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_sample_start_
      -- 
    req_3277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(329), ack => WPIPE_ConvTranspose_output_pipe_1534_inst_req_0); -- 
    convTranspose_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(309) & convTranspose_CP_772_elements(328);
      gj_convTranspose_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  transition  input  output  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (6) 
      -- CP-element group 330: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Update/req
      -- CP-element group 330: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Sample/ack
      -- CP-element group 330: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_update_start_
      -- CP-element group 330: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_sample_completed_
      -- 
    ack_3278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1534_inst_ack_0, ack => convTranspose_CP_772_elements(330)); -- 
    req_3282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(330), ack => WPIPE_ConvTranspose_output_pipe_1534_inst_req_1); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Update/ack
      -- CP-element group 331: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1534_update_completed_
      -- 
    ack_3283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1534_inst_ack_1, ack => convTranspose_CP_772_elements(331)); -- 
    -- CP-element group 332:  join  transition  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	307 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Sample/req
      -- CP-element group 332: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Sample/$entry
      -- 
    req_3291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(332), ack => WPIPE_ConvTranspose_output_pipe_1537_inst_req_0); -- 
    convTranspose_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(307) & convTranspose_CP_772_elements(331);
      gj_convTranspose_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_update_start_
      -- CP-element group 333: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Update/req
      -- CP-element group 333: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Sample/ack
      -- 
    ack_3292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1537_inst_ack_0, ack => convTranspose_CP_772_elements(333)); -- 
    req_3296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(333), ack => WPIPE_ConvTranspose_output_pipe_1537_inst_req_1); -- 
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1537_Update/$exit
      -- 
    ack_3297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1537_inst_ack_1, ack => convTranspose_CP_772_elements(334)); -- 
    -- CP-element group 335:  join  transition  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	305 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Sample/req
      -- CP-element group 335: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_sample_start_
      -- 
    req_3305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(335), ack => WPIPE_ConvTranspose_output_pipe_1540_inst_req_0); -- 
    convTranspose_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(305) & convTranspose_CP_772_elements(334);
      gj_convTranspose_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_sample_completed_
      -- CP-element group 336: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Sample/$exit
      -- CP-element group 336: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_update_start_
      -- CP-element group 336: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Update/req
      -- CP-element group 336: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Sample/ack
      -- 
    ack_3306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1540_inst_ack_0, ack => convTranspose_CP_772_elements(336)); -- 
    req_3310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(336), ack => WPIPE_ConvTranspose_output_pipe_1540_inst_req_1); -- 
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Update/ack
      -- CP-element group 337: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1540_Update/$exit
      -- 
    ack_3311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1540_inst_ack_1, ack => convTranspose_CP_772_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	303 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Sample/req
      -- CP-element group 338: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_sample_start_
      -- 
    req_3319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(338), ack => WPIPE_ConvTranspose_output_pipe_1543_inst_req_0); -- 
    convTranspose_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(303) & convTranspose_CP_772_elements(337);
      gj_convTranspose_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_update_start_
      -- CP-element group 339: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Update/req
      -- 
    ack_3320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1543_inst_ack_0, ack => convTranspose_CP_772_elements(339)); -- 
    req_3324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(339), ack => WPIPE_ConvTranspose_output_pipe_1543_inst_req_1); -- 
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/WPIPE_ConvTranspose_output_pipe_1543_Update/ack
      -- 
    ack_3325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1543_inst_ack_1, ack => convTranspose_CP_772_elements(340)); -- 
    -- CP-element group 341:  branch  join  transition  place  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	296 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: 	343 
    -- CP-element group 341:  members (10) 
      -- CP-element group 341: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556__exit__
      -- CP-element group 341: 	 branch_block_stmt_312/if_stmt_1557__entry__
      -- CP-element group 341: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/$exit
      -- CP-element group 341: 	 branch_block_stmt_312/if_stmt_1557_dead_link/$entry
      -- CP-element group 341: 	 branch_block_stmt_312/if_stmt_1557_eval_test/$entry
      -- CP-element group 341: 	 branch_block_stmt_312/if_stmt_1557_eval_test/$exit
      -- CP-element group 341: 	 branch_block_stmt_312/if_stmt_1557_eval_test/branch_req
      -- CP-element group 341: 	 branch_block_stmt_312/R_exitcond8_1558_place
      -- CP-element group 341: 	 branch_block_stmt_312/if_stmt_1557_if_link/$entry
      -- CP-element group 341: 	 branch_block_stmt_312/if_stmt_1557_else_link/$entry
      -- 
    branch_req_3333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(341), ack => if_stmt_1557_branch_req_0); -- 
    convTranspose_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(296) & convTranspose_CP_772_elements(340);
      gj_convTranspose_cp_element_group_341 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  merge  transition  place  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	371 
    -- CP-element group 342:  members (13) 
      -- CP-element group 342: 	 branch_block_stmt_312/merge_stmt_1563__exit__
      -- CP-element group 342: 	 branch_block_stmt_312/forx_xend417x_xloopexit_forx_xend417
      -- CP-element group 342: 	 branch_block_stmt_312/if_stmt_1557_if_link/$exit
      -- CP-element group 342: 	 branch_block_stmt_312/if_stmt_1557_if_link/if_choice_transition
      -- CP-element group 342: 	 branch_block_stmt_312/forx_xbody345_forx_xend417x_xloopexit
      -- CP-element group 342: 	 branch_block_stmt_312/forx_xbody345_forx_xend417x_xloopexit_PhiReq/$entry
      -- CP-element group 342: 	 branch_block_stmt_312/forx_xbody345_forx_xend417x_xloopexit_PhiReq/$exit
      -- CP-element group 342: 	 branch_block_stmt_312/merge_stmt_1563_PhiReqMerge
      -- CP-element group 342: 	 branch_block_stmt_312/merge_stmt_1563_PhiAck/$entry
      -- CP-element group 342: 	 branch_block_stmt_312/merge_stmt_1563_PhiAck/$exit
      -- CP-element group 342: 	 branch_block_stmt_312/merge_stmt_1563_PhiAck/dummy
      -- CP-element group 342: 	 branch_block_stmt_312/forx_xend417x_xloopexit_forx_xend417_PhiReq/$entry
      -- CP-element group 342: 	 branch_block_stmt_312/forx_xend417x_xloopexit_forx_xend417_PhiReq/$exit
      -- 
    if_choice_transition_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1557_branch_ack_1, ack => convTranspose_CP_772_elements(342)); -- 
    -- CP-element group 343:  fork  transition  place  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	341 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	366 
    -- CP-element group 343: 	367 
    -- CP-element group 343:  members (12) 
      -- CP-element group 343: 	 branch_block_stmt_312/if_stmt_1557_else_link/$exit
      -- CP-element group 343: 	 branch_block_stmt_312/if_stmt_1557_else_link/else_choice_transition
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/$entry
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/$entry
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$entry
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/$entry
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/$entry
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Sample/rr
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1557_branch_ack_0, ack => convTranspose_CP_772_elements(343)); -- 
    rr_3617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(343), ack => type_cast_1433_inst_req_0); -- 
    cr_3622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(343), ack => type_cast_1433_inst_req_1); -- 
    -- CP-element group 344:  merge  branch  transition  place  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	164 
    -- CP-element group 344: 	114 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	115 
    -- CP-element group 344: 	116 
    -- CP-element group 344:  members (17) 
      -- CP-element group 344: 	 branch_block_stmt_312/merge_stmt_672__exit__
      -- CP-element group 344: 	 branch_block_stmt_312/assign_stmt_678__entry__
      -- CP-element group 344: 	 branch_block_stmt_312/assign_stmt_678__exit__
      -- CP-element group 344: 	 branch_block_stmt_312/if_stmt_679__entry__
      -- CP-element group 344: 	 branch_block_stmt_312/assign_stmt_678/$entry
      -- CP-element group 344: 	 branch_block_stmt_312/assign_stmt_678/$exit
      -- CP-element group 344: 	 branch_block_stmt_312/if_stmt_679_dead_link/$entry
      -- CP-element group 344: 	 branch_block_stmt_312/if_stmt_679_eval_test/$entry
      -- CP-element group 344: 	 branch_block_stmt_312/if_stmt_679_eval_test/$exit
      -- CP-element group 344: 	 branch_block_stmt_312/if_stmt_679_eval_test/branch_req
      -- CP-element group 344: 	 branch_block_stmt_312/R_cmp180426_680_place
      -- CP-element group 344: 	 branch_block_stmt_312/if_stmt_679_if_link/$entry
      -- CP-element group 344: 	 branch_block_stmt_312/if_stmt_679_else_link/$entry
      -- CP-element group 344: 	 branch_block_stmt_312/merge_stmt_672_PhiReqMerge
      -- CP-element group 344: 	 branch_block_stmt_312/merge_stmt_672_PhiAck/$entry
      -- CP-element group 344: 	 branch_block_stmt_312/merge_stmt_672_PhiAck/$exit
      -- CP-element group 344: 	 branch_block_stmt_312/merge_stmt_672_PhiAck/dummy
      -- 
    branch_req_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(344), ack => if_stmt_679_branch_req_0); -- 
    convTranspose_CP_772_elements(344) <= OrReduce(convTranspose_CP_772_elements(164) & convTranspose_CP_772_elements(114));
    -- CP-element group 345:  transition  output  delay-element  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	123 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	349 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/$exit
      -- CP-element group 345: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/phi_stmt_729/$exit
      -- CP-element group 345: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/$exit
      -- CP-element group 345: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_733_konst_delay_trans
      -- CP-element group 345: 	 branch_block_stmt_312/bbx_xnph432_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_req
      -- 
    phi_stmt_729_req_3390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_729_req_3390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(345), ack => phi_stmt_729_req_0); -- 
    -- Element group convTranspose_CP_772_elements(345) is a control-delay.
    cp_element_345_delay: control_delay_element  generic map(name => " 345_delay", delay_value => 1)  port map(req => convTranspose_CP_772_elements(123), ack => convTranspose_CP_772_elements(345), clk => clk, reset =>reset);
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	165 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Sample/ra
      -- 
    ra_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_0, ack => convTranspose_CP_772_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	165 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (2) 
      -- CP-element group 347: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/Update/ca
      -- 
    ca_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_1, ack => convTranspose_CP_772_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (6) 
      -- CP-element group 348: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 348: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/$exit
      -- CP-element group 348: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/$exit
      -- CP-element group 348: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/$exit
      -- CP-element group 348: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_sources/type_cast_735/SplitProtocol/$exit
      -- CP-element group 348: 	 branch_block_stmt_312/forx_xbody_forx_xbody_PhiReq/phi_stmt_729/phi_stmt_729_req
      -- 
    phi_stmt_729_req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_729_req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(348), ack => phi_stmt_729_req_1); -- 
    convTranspose_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(346) & convTranspose_CP_772_elements(347);
      gj_convTranspose_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  merge  transition  place  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	345 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (2) 
      -- CP-element group 349: 	 branch_block_stmt_312/merge_stmt_728_PhiReqMerge
      -- CP-element group 349: 	 branch_block_stmt_312/merge_stmt_728_PhiAck/$entry
      -- 
    convTranspose_CP_772_elements(349) <= OrReduce(convTranspose_CP_772_elements(345) & convTranspose_CP_772_elements(348));
    -- CP-element group 350:  fork  transition  place  input  output  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	155 
    -- CP-element group 350: 	159 
    -- CP-element group 350: 	162 
    -- CP-element group 350: 	124 
    -- CP-element group 350: 	125 
    -- CP-element group 350: 	127 
    -- CP-element group 350: 	128 
    -- CP-element group 350: 	131 
    -- CP-element group 350: 	135 
    -- CP-element group 350: 	139 
    -- CP-element group 350: 	143 
    -- CP-element group 350: 	147 
    -- CP-element group 350: 	151 
    -- CP-element group 350:  members (56) 
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/word_access_complete/word_0/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/word_access_complete/word_0/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/word_access_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/merge_stmt_728__exit__
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893__entry__
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/ptr_deref_880_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_836_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_872_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_resized_2
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_scaled_2
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_computed_2
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_resize_2/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_resize_2/$exit
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_resize_2/index_resize_req
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_resize_2/index_resize_ack
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_scale_2/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_scale_2/$exit
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_scale_2/scale_rename_req
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_index_scale_2/scale_rename_ack
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_update_start
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Sample/req
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/array_obj_ref_743_final_index_sum_regn_Update/req
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/addr_of_744_complete/req
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_sample_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/RPIPE_ConvTranspose_input_pipe_747_Sample/rr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_751_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_764_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_854_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_782_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_818_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_312/assign_stmt_745_to_assign_stmt_893/type_cast_800_update_start_
      -- CP-element group 350: 	 branch_block_stmt_312/merge_stmt_728_PhiAck/$exit
      -- CP-element group 350: 	 branch_block_stmt_312/merge_stmt_728_PhiAck/phi_stmt_729_ack
      -- 
    phi_stmt_729_ack_3421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_729_ack_0, ack => convTranspose_CP_772_elements(350)); -- 
    cr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => ptr_deref_880_store_0_req_1); -- 
    cr_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_800_inst_req_1); -- 
    cr_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_836_inst_req_1); -- 
    cr_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_872_inst_req_1); -- 
    req_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => array_obj_ref_743_index_offset_req_0); -- 
    req_1723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => array_obj_ref_743_index_offset_req_1); -- 
    req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => addr_of_744_final_reg_req_1); -- 
    rr_1747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => RPIPE_ConvTranspose_input_pipe_747_inst_req_0); -- 
    cr_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_751_inst_req_1); -- 
    cr_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_854_inst_req_1); -- 
    cr_1794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_764_inst_req_1); -- 
    cr_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_818_inst_req_1); -- 
    cr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(350), ack => type_cast_782_inst_req_1); -- 
    -- CP-element group 351:  transition  output  delay-element  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	170 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	355 
    -- CP-element group 351:  members (5) 
      -- CP-element group 351: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/$exit
      -- CP-element group 351: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/phi_stmt_945/$exit
      -- CP-element group 351: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/$exit
      -- CP-element group 351: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_951_konst_delay_trans
      -- CP-element group 351: 	 branch_block_stmt_312/bbx_xnph428_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_req
      -- 
    phi_stmt_945_req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_945_req_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(351), ack => phi_stmt_945_req_1); -- 
    -- Element group convTranspose_CP_772_elements(351) is a control-delay.
    cp_element_351_delay: control_delay_element  generic map(name => " 351_delay", delay_value => 1)  port map(req => convTranspose_CP_772_elements(170), ack => convTranspose_CP_772_elements(351), clk => clk, reset =>reset);
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	212 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	354 
    -- CP-element group 352:  members (2) 
      -- CP-element group 352: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/ra
      -- 
    ra_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_948_inst_ack_0, ack => convTranspose_CP_772_elements(352)); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	212 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (2) 
      -- CP-element group 353: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/ca
      -- 
    ca_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_948_inst_ack_1, ack => convTranspose_CP_772_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	352 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (6) 
      -- CP-element group 354: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/$exit
      -- CP-element group 354: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/$exit
      -- CP-element group 354: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/$exit
      -- CP-element group 354: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/$exit
      -- CP-element group 354: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/$exit
      -- CP-element group 354: 	 branch_block_stmt_312/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_945/phi_stmt_945_req
      -- 
    phi_stmt_945_req_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_945_req_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(354), ack => phi_stmt_945_req_0); -- 
    convTranspose_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(352) & convTranspose_CP_772_elements(353);
      gj_convTranspose_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  merge  transition  place  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	351 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (2) 
      -- CP-element group 355: 	 branch_block_stmt_312/merge_stmt_944_PhiReqMerge
      -- CP-element group 355: 	 branch_block_stmt_312/merge_stmt_944_PhiAck/$entry
      -- 
    convTranspose_CP_772_elements(355) <= OrReduce(convTranspose_CP_772_elements(351) & convTranspose_CP_772_elements(354));
    -- CP-element group 356:  fork  transition  place  input  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	209 
    -- CP-element group 356: 	198 
    -- CP-element group 356: 	202 
    -- CP-element group 356: 	206 
    -- CP-element group 356: 	171 
    -- CP-element group 356: 	172 
    -- CP-element group 356: 	174 
    -- CP-element group 356: 	175 
    -- CP-element group 356: 	178 
    -- CP-element group 356: 	182 
    -- CP-element group 356: 	186 
    -- CP-element group 356: 	190 
    -- CP-element group 356: 	194 
    -- CP-element group 356:  members (56) 
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_complete/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_complete/req
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Update/req
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/merge_stmt_944__exit__
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109__entry__
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Sample/req
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_final_index_sum_regn_update_start
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_998_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_scale_2/scale_rename_ack
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_980_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_scale_2/scale_rename_req
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_scale_2/$exit
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_scale_2/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_resize_2/index_resize_ack
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_resize_2/index_resize_req
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_resize_2/$exit
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_resize_2/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_computed_2
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_scaled_2
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/array_obj_ref_959_index_resized_2
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/addr_of_960_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1052_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1034_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1070_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_967_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Sample/rr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/RPIPE_ConvTranspose_input_pipe_963_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1016_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/type_cast_1088_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_update_start_
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/word_access_complete/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/word_access_complete/word_0/$entry
      -- CP-element group 356: 	 branch_block_stmt_312/assign_stmt_961_to_assign_stmt_1109/ptr_deref_1096_Update/word_access_complete/word_0/cr
      -- CP-element group 356: 	 branch_block_stmt_312/merge_stmt_944_PhiAck/$exit
      -- CP-element group 356: 	 branch_block_stmt_312/merge_stmt_944_PhiAck/phi_stmt_945_ack
      -- 
    phi_stmt_945_ack_3475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_945_ack_0, ack => convTranspose_CP_772_elements(356)); -- 
    cr_2195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_998_inst_req_1); -- 
    cr_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_1016_inst_req_1); -- 
    cr_2251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_1034_inst_req_1); -- 
    req_2111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => addr_of_960_final_reg_req_1); -- 
    cr_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_980_inst_req_1); -- 
    req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => array_obj_ref_959_index_offset_req_1); -- 
    req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => array_obj_ref_959_index_offset_req_0); -- 
    cr_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_1052_inst_req_1); -- 
    cr_2139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_967_inst_req_1); -- 
    cr_2307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_1070_inst_req_1); -- 
    rr_2120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => RPIPE_ConvTranspose_input_pipe_963_inst_req_0); -- 
    cr_2335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => type_cast_1088_inst_req_1); -- 
    cr_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(356), ack => ptr_deref_1096_store_0_req_1); -- 
    -- CP-element group 357:  merge  fork  transition  place  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	211 
    -- CP-element group 357: 	116 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	213 
    -- CP-element group 357: 	214 
    -- CP-element group 357: 	215 
    -- CP-element group 357: 	216 
    -- CP-element group 357: 	217 
    -- CP-element group 357: 	218 
    -- CP-element group 357:  members (25) 
      -- CP-element group 357: 	 branch_block_stmt_312/merge_stmt_1118__exit__
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146__entry__
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_update_start_
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Sample/rr
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1121_Update/cr
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_update_start_
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Sample/rr
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1125_Update/cr
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_update_start_
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Sample/rr
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/assign_stmt_1122_to_assign_stmt_1146/type_cast_1129_Update/cr
      -- CP-element group 357: 	 branch_block_stmt_312/merge_stmt_1118_PhiReqMerge
      -- CP-element group 357: 	 branch_block_stmt_312/merge_stmt_1118_PhiAck/$entry
      -- CP-element group 357: 	 branch_block_stmt_312/merge_stmt_1118_PhiAck/$exit
      -- CP-element group 357: 	 branch_block_stmt_312/merge_stmt_1118_PhiAck/dummy
      -- 
    rr_2416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(357), ack => type_cast_1121_inst_req_0); -- 
    cr_2421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(357), ack => type_cast_1121_inst_req_1); -- 
    rr_2430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(357), ack => type_cast_1125_inst_req_0); -- 
    cr_2435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(357), ack => type_cast_1125_inst_req_1); -- 
    rr_2444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(357), ack => type_cast_1129_inst_req_0); -- 
    cr_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(357), ack => type_cast_1129_inst_req_1); -- 
    convTranspose_CP_772_elements(357) <= OrReduce(convTranspose_CP_772_elements(211) & convTranspose_CP_772_elements(116));
    -- CP-element group 358:  transition  output  delay-element  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	228 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	362 
    -- CP-element group 358:  members (5) 
      -- CP-element group 358: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/$exit
      -- CP-element group 358: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/phi_stmt_1197/$exit
      -- CP-element group 358: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/$exit
      -- CP-element group 358: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1201_konst_delay_trans
      -- CP-element group 358: 	 branch_block_stmt_312/bbx_xnph424_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_req
      -- 
    phi_stmt_1197_req_3521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1197_req_3521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(358), ack => phi_stmt_1197_req_0); -- 
    -- Element group convTranspose_CP_772_elements(358) is a control-delay.
    cp_element_358_delay: control_delay_element  generic map(name => " 358_delay", delay_value => 1)  port map(req => convTranspose_CP_772_elements(228), ack => convTranspose_CP_772_elements(358), clk => clk, reset =>reset);
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	237 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (2) 
      -- CP-element group 359: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Sample/ra
      -- 
    ra_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_0, ack => convTranspose_CP_772_elements(359)); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	237 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (2) 
      -- CP-element group 360: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/Update/ca
      -- 
    ca_3546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_1, ack => convTranspose_CP_772_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/$exit
      -- CP-element group 361: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/$exit
      -- CP-element group 361: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/$exit
      -- CP-element group 361: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/$exit
      -- CP-element group 361: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_sources/type_cast_1203/SplitProtocol/$exit
      -- CP-element group 361: 	 branch_block_stmt_312/forx_xbody251_forx_xbody251_PhiReq/phi_stmt_1197/phi_stmt_1197_req
      -- 
    phi_stmt_1197_req_3547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1197_req_3547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(361), ack => phi_stmt_1197_req_1); -- 
    convTranspose_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(359) & convTranspose_CP_772_elements(360);
      gj_convTranspose_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  merge  transition  place  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	358 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_312/merge_stmt_1196_PhiReqMerge
      -- CP-element group 362: 	 branch_block_stmt_312/merge_stmt_1196_PhiAck/$entry
      -- 
    convTranspose_CP_772_elements(362) <= OrReduce(convTranspose_CP_772_elements(358) & convTranspose_CP_772_elements(361));
    -- CP-element group 363:  fork  transition  place  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	229 
    -- CP-element group 363: 	230 
    -- CP-element group 363: 	232 
    -- CP-element group 363: 	234 
    -- CP-element group 363:  members (29) 
      -- CP-element group 363: 	 branch_block_stmt_312/merge_stmt_1196__exit__
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229__entry__
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_update_start_
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_resized_2
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_scaled_2
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_computed_2
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_resize_2/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_resize_2/$exit
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_resize_2/index_resize_req
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_resize_2/index_resize_ack
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_scale_2/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_scale_2/$exit
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_scale_2/scale_rename_req
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_index_scale_2/scale_rename_ack
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_update_start
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Sample/req
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/array_obj_ref_1211_final_index_sum_regn_Update/req
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_complete/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/addr_of_1212_complete/req
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_update_start_
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/word_access_complete/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/word_access_complete/word_0/$entry
      -- CP-element group 363: 	 branch_block_stmt_312/assign_stmt_1213_to_assign_stmt_1229/ptr_deref_1215_Update/word_access_complete/word_0/cr
      -- CP-element group 363: 	 branch_block_stmt_312/merge_stmt_1196_PhiAck/$exit
      -- CP-element group 363: 	 branch_block_stmt_312/merge_stmt_1196_PhiAck/phi_stmt_1197_ack
      -- 
    phi_stmt_1197_ack_3552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1197_ack_0, ack => convTranspose_CP_772_elements(363)); -- 
    req_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(363), ack => array_obj_ref_1211_index_offset_req_0); -- 
    req_2547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(363), ack => array_obj_ref_1211_index_offset_req_1); -- 
    req_2562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(363), ack => addr_of_1212_final_reg_req_1); -- 
    cr_2612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(363), ack => ptr_deref_1215_store_0_req_1); -- 
    -- CP-element group 364:  merge  fork  transition  place  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	221 
    -- CP-element group 364: 	236 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	238 
    -- CP-element group 364: 	239 
    -- CP-element group 364: 	241 
    -- CP-element group 364:  members (16) 
      -- CP-element group 364: 	 branch_block_stmt_312/merge_stmt_1238__exit__
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247__entry__
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/$entry
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_sample_start_
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_update_start_
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Sample/$entry
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Sample/crr
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Update/$entry
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/call_stmt_1241_Update/ccr
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_update_start_
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Update/$entry
      -- CP-element group 364: 	 branch_block_stmt_312/call_stmt_1241_to_assign_stmt_1247/type_cast_1246_Update/cr
      -- CP-element group 364: 	 branch_block_stmt_312/merge_stmt_1238_PhiReqMerge
      -- CP-element group 364: 	 branch_block_stmt_312/merge_stmt_1238_PhiAck/$entry
      -- CP-element group 364: 	 branch_block_stmt_312/merge_stmt_1238_PhiAck/$exit
      -- CP-element group 364: 	 branch_block_stmt_312/merge_stmt_1238_PhiAck/dummy
      -- 
    crr_2643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(364), ack => call_stmt_1241_call_req_0); -- 
    ccr_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(364), ack => call_stmt_1241_call_req_1); -- 
    cr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(364), ack => type_cast_1246_inst_req_1); -- 
    convTranspose_CP_772_elements(364) <= OrReduce(convTranspose_CP_772_elements(221) & convTranspose_CP_772_elements(236));
    -- CP-element group 365:  transition  output  delay-element  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	295 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	369 
    -- CP-element group 365:  members (5) 
      -- CP-element group 365: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/$exit
      -- CP-element group 365: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/phi_stmt_1427/$exit
      -- CP-element group 365: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$exit
      -- CP-element group 365: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1431_konst_delay_trans
      -- CP-element group 365: 	 branch_block_stmt_312/bbx_xnph_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_req
      -- 
    phi_stmt_1427_req_3598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1427_req_3598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(365), ack => phi_stmt_1427_req_0); -- 
    -- Element group convTranspose_CP_772_elements(365) is a control-delay.
    cp_element_365_delay: control_delay_element  generic map(name => " 365_delay", delay_value => 1)  port map(req => convTranspose_CP_772_elements(295), ack => convTranspose_CP_772_elements(365), clk => clk, reset =>reset);
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	343 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (2) 
      -- CP-element group 366: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Sample/ra
      -- 
    ra_3618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1433_inst_ack_0, ack => convTranspose_CP_772_elements(366)); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	343 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/Update/ca
      -- 
    ca_3623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1433_inst_ack_1, ack => convTranspose_CP_772_elements(367)); -- 
    -- CP-element group 368:  join  transition  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/$exit
      -- CP-element group 368: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/$exit
      -- CP-element group 368: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$exit
      -- CP-element group 368: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/$exit
      -- CP-element group 368: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433/SplitProtocol/$exit
      -- CP-element group 368: 	 branch_block_stmt_312/forx_xbody345_forx_xbody345_PhiReq/phi_stmt_1427/phi_stmt_1427_req
      -- 
    phi_stmt_1427_req_3624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1427_req_3624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(368), ack => phi_stmt_1427_req_1); -- 
    convTranspose_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_772_elements(366) & convTranspose_CP_772_elements(367);
      gj_convTranspose_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_772_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  merge  transition  place  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	365 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_312/merge_stmt_1426_PhiReqMerge
      -- CP-element group 369: 	 branch_block_stmt_312/merge_stmt_1426_PhiAck/$entry
      -- 
    convTranspose_CP_772_elements(369) <= OrReduce(convTranspose_CP_772_elements(365) & convTranspose_CP_772_elements(368));
    -- CP-element group 370:  fork  transition  place  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	296 
    -- CP-element group 370: 	297 
    -- CP-element group 370: 	299 
    -- CP-element group 370: 	301 
    -- CP-element group 370: 	303 
    -- CP-element group 370: 	305 
    -- CP-element group 370: 	307 
    -- CP-element group 370: 	309 
    -- CP-element group 370: 	311 
    -- CP-element group 370: 	313 
    -- CP-element group 370: 	315 
    -- CP-element group 370: 	317 
    -- CP-element group 370:  members (53) 
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/merge_stmt_1426__exit__
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556__entry__
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1500_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_resized_2
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1480_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1470_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_complete/req
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1460_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/addr_of_1442_complete/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1490_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1510_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Update/req
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1450_update_start_
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Sample/req
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_final_index_sum_regn_update_start
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_scale_2/scale_rename_ack
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_scale_2/scale_rename_req
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/word_access_complete/word_0/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/word_access_complete/word_0/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_scale_2/$exit
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_scale_2/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/word_access_complete/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_resize_2/index_resize_ack
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_resize_2/index_resize_req
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/ptr_deref_1446_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_resize_2/$exit
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_resize_2/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_computed_2
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/type_cast_1520_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_312/assign_stmt_1443_to_assign_stmt_1556/array_obj_ref_1441_index_scaled_2
      -- CP-element group 370: 	 branch_block_stmt_312/merge_stmt_1426_PhiAck/$exit
      -- CP-element group 370: 	 branch_block_stmt_312/merge_stmt_1426_PhiAck/phi_stmt_1427_ack
      -- 
    phi_stmt_1427_ack_3629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1427_ack_0, ack => convTranspose_CP_772_elements(370)); -- 
    cr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1500_inst_req_1); -- 
    cr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1480_inst_req_1); -- 
    cr_3142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1470_inst_req_1); -- 
    cr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1490_inst_req_1); -- 
    cr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1510_inst_req_1); -- 
    cr_3128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1460_inst_req_1); -- 
    req_3050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => addr_of_1442_final_reg_req_1); -- 
    cr_3114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1450_inst_req_1); -- 
    req_3035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => array_obj_ref_1441_index_offset_req_1); -- 
    req_3030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => array_obj_ref_1441_index_offset_req_0); -- 
    cr_3095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => ptr_deref_1446_load_0_req_1); -- 
    cr_3212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_772_elements(370), ack => type_cast_1520_inst_req_1); -- 
    -- CP-element group 371:  merge  transition  place  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	288 
    -- CP-element group 371: 	342 
    -- CP-element group 371: successors 
    -- CP-element group 371:  members (16) 
      -- CP-element group 371: 	 $exit
      -- CP-element group 371: 	 branch_block_stmt_312/$exit
      -- CP-element group 371: 	 branch_block_stmt_312/branch_block_stmt_312__exit__
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1565__exit__
      -- CP-element group 371: 	 branch_block_stmt_312/return__
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1567__exit__
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1565_PhiReqMerge
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1565_PhiAck/$entry
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1565_PhiAck/$exit
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1565_PhiAck/dummy
      -- CP-element group 371: 	 branch_block_stmt_312/return___PhiReq/$entry
      -- CP-element group 371: 	 branch_block_stmt_312/return___PhiReq/$exit
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1567_PhiReqMerge
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1567_PhiAck/$entry
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1567_PhiAck/$exit
      -- CP-element group 371: 	 branch_block_stmt_312/merge_stmt_1567_PhiAck/dummy
      -- 
    convTranspose_CP_772_elements(371) <= OrReduce(convTranspose_CP_772_elements(288) & convTranspose_CP_772_elements(342));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_ix_x0431_742_resized : std_logic_vector(15 downto 0);
    signal R_ix_x0431_742_scaled : std_logic_vector(15 downto 0);
    signal R_ix_x1427_958_resized : std_logic_vector(15 downto 0);
    signal R_ix_x1427_958_scaled : std_logic_vector(15 downto 0);
    signal R_ix_x2423_1210_resized : std_logic_vector(15 downto 0);
    signal R_ix_x2423_1210_scaled : std_logic_vector(15 downto 0);
    signal R_ix_x3420_1440_resized : std_logic_vector(15 downto 0);
    signal R_ix_x3420_1440_scaled : std_logic_vector(15 downto 0);
    signal add104_607 : std_logic_vector(15 downto 0);
    signal add113_632 : std_logic_vector(15 downto 0);
    signal add122_657 : std_logic_vector(15 downto 0);
    signal add12_362 : std_logic_vector(15 downto 0);
    signal add136_770 : std_logic_vector(63 downto 0);
    signal add142_788 : std_logic_vector(63 downto 0);
    signal add148_806 : std_logic_vector(63 downto 0);
    signal add154_824 : std_logic_vector(63 downto 0);
    signal add160_842 : std_logic_vector(63 downto 0);
    signal add166_860 : std_logic_vector(63 downto 0);
    signal add172_878 : std_logic_vector(63 downto 0);
    signal add192_986 : std_logic_vector(63 downto 0);
    signal add198_1004 : std_logic_vector(63 downto 0);
    signal add204_1022 : std_logic_vector(63 downto 0);
    signal add210_1040 : std_logic_vector(63 downto 0);
    signal add216_1058 : std_logic_vector(63 downto 0);
    signal add21_387 : std_logic_vector(15 downto 0);
    signal add222_1076 : std_logic_vector(63 downto 0);
    signal add228_1094 : std_logic_vector(63 downto 0);
    signal add30_412 : std_logic_vector(31 downto 0);
    signal add39_437 : std_logic_vector(15 downto 0);
    signal add48_462 : std_logic_vector(15 downto 0);
    signal add57_487 : std_logic_vector(31 downto 0);
    signal add86_557 : std_logic_vector(15 downto 0);
    signal add95_582 : std_logic_vector(15 downto 0);
    signal add_337 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1211_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1211_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1211_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1211_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1211_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1211_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1211_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1441_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1441_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1441_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1441_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1441_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1441_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1441_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_743_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_743_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_743_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_743_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_743_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_743_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_743_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_959_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_959_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_959_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_959_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_959_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_959_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_959_root_address : std_logic_vector(15 downto 0);
    signal arrayidx231_961 : std_logic_vector(31 downto 0);
    signal arrayidx253_1213 : std_logic_vector(31 downto 0);
    signal arrayidx349_1443 : std_logic_vector(31 downto 0);
    signal arrayidx_745 : std_logic_vector(31 downto 0);
    signal call102_598 : std_logic_vector(7 downto 0);
    signal call106_610 : std_logic_vector(7 downto 0);
    signal call10_353 : std_logic_vector(7 downto 0);
    signal call111_623 : std_logic_vector(7 downto 0);
    signal call115_635 : std_logic_vector(7 downto 0);
    signal call120_648 : std_logic_vector(7 downto 0);
    signal call129_748 : std_logic_vector(7 downto 0);
    signal call133_761 : std_logic_vector(7 downto 0);
    signal call139_779 : std_logic_vector(7 downto 0);
    signal call145_797 : std_logic_vector(7 downto 0);
    signal call14_365 : std_logic_vector(7 downto 0);
    signal call151_815 : std_logic_vector(7 downto 0);
    signal call157_833 : std_logic_vector(7 downto 0);
    signal call163_851 : std_logic_vector(7 downto 0);
    signal call169_869 : std_logic_vector(7 downto 0);
    signal call185_964 : std_logic_vector(7 downto 0);
    signal call189_977 : std_logic_vector(7 downto 0);
    signal call195_995 : std_logic_vector(7 downto 0);
    signal call19_378 : std_logic_vector(7 downto 0);
    signal call201_1013 : std_logic_vector(7 downto 0);
    signal call207_1031 : std_logic_vector(7 downto 0);
    signal call213_1049 : std_logic_vector(7 downto 0);
    signal call219_1067 : std_logic_vector(7 downto 0);
    signal call225_1085 : std_logic_vector(7 downto 0);
    signal call23_390 : std_logic_vector(7 downto 0);
    signal call259_1241 : std_logic_vector(63 downto 0);
    signal call272_1266 : std_logic_vector(63 downto 0);
    signal call28_403 : std_logic_vector(7 downto 0);
    signal call2_328 : std_logic_vector(7 downto 0);
    signal call32_415 : std_logic_vector(7 downto 0);
    signal call37_428 : std_logic_vector(7 downto 0);
    signal call41_440 : std_logic_vector(7 downto 0);
    signal call46_453 : std_logic_vector(7 downto 0);
    signal call50_465 : std_logic_vector(7 downto 0);
    signal call55_478 : std_logic_vector(7 downto 0);
    signal call5_340 : std_logic_vector(7 downto 0);
    signal call79_535 : std_logic_vector(7 downto 0);
    signal call84_548 : std_logic_vector(7 downto 0);
    signal call88_560 : std_logic_vector(7 downto 0);
    signal call93_573 : std_logic_vector(7 downto 0);
    signal call97_585 : std_logic_vector(7 downto 0);
    signal call_315 : std_logic_vector(7 downto 0);
    signal cmp180426_678 : std_logic_vector(0 downto 0);
    signal cmp249422_1146 : std_logic_vector(0 downto 0);
    signal cmp430_663 : std_logic_vector(0 downto 0);
    signal conv100_589 : std_logic_vector(15 downto 0);
    signal conv103_602 : std_logic_vector(15 downto 0);
    signal conv109_614 : std_logic_vector(15 downto 0);
    signal conv112_627 : std_logic_vector(15 downto 0);
    signal conv118_639 : std_logic_vector(15 downto 0);
    signal conv11_357 : std_logic_vector(15 downto 0);
    signal conv121_652 : std_logic_vector(15 downto 0);
    signal conv130_752 : std_logic_vector(63 downto 0);
    signal conv135_765 : std_logic_vector(63 downto 0);
    signal conv141_783 : std_logic_vector(63 downto 0);
    signal conv147_801 : std_logic_vector(63 downto 0);
    signal conv153_819 : std_logic_vector(63 downto 0);
    signal conv159_837 : std_logic_vector(63 downto 0);
    signal conv165_855 : std_logic_vector(63 downto 0);
    signal conv171_873 : std_logic_vector(63 downto 0);
    signal conv17_369 : std_logic_vector(15 downto 0);
    signal conv186_968 : std_logic_vector(63 downto 0);
    signal conv191_981 : std_logic_vector(63 downto 0);
    signal conv197_999 : std_logic_vector(63 downto 0);
    signal conv1_319 : std_logic_vector(15 downto 0);
    signal conv203_1017 : std_logic_vector(63 downto 0);
    signal conv209_1035 : std_logic_vector(63 downto 0);
    signal conv20_382 : std_logic_vector(15 downto 0);
    signal conv215_1053 : std_logic_vector(63 downto 0);
    signal conv221_1071 : std_logic_vector(63 downto 0);
    signal conv227_1089 : std_logic_vector(63 downto 0);
    signal conv238_1122 : std_logic_vector(31 downto 0);
    signal conv240_1126 : std_logic_vector(31 downto 0);
    signal conv243_1130 : std_logic_vector(31 downto 0);
    signal conv260_1247 : std_logic_vector(63 downto 0);
    signal conv26_394 : std_logic_vector(31 downto 0);
    signal conv273_1271 : std_logic_vector(63 downto 0);
    signal conv279_1281 : std_logic_vector(7 downto 0);
    signal conv285_1291 : std_logic_vector(7 downto 0);
    signal conv291_1301 : std_logic_vector(7 downto 0);
    signal conv297_1311 : std_logic_vector(7 downto 0);
    signal conv29_407 : std_logic_vector(31 downto 0);
    signal conv303_1321 : std_logic_vector(7 downto 0);
    signal conv309_1331 : std_logic_vector(7 downto 0);
    signal conv315_1341 : std_logic_vector(7 downto 0);
    signal conv321_1351 : std_logic_vector(7 downto 0);
    signal conv354_1451 : std_logic_vector(7 downto 0);
    signal conv35_419 : std_logic_vector(15 downto 0);
    signal conv360_1461 : std_logic_vector(7 downto 0);
    signal conv366_1471 : std_logic_vector(7 downto 0);
    signal conv372_1481 : std_logic_vector(7 downto 0);
    signal conv378_1491 : std_logic_vector(7 downto 0);
    signal conv384_1501 : std_logic_vector(7 downto 0);
    signal conv38_432 : std_logic_vector(15 downto 0);
    signal conv390_1511 : std_logic_vector(7 downto 0);
    signal conv396_1521 : std_logic_vector(7 downto 0);
    signal conv3_332 : std_logic_vector(15 downto 0);
    signal conv44_444 : std_logic_vector(15 downto 0);
    signal conv47_457 : std_logic_vector(15 downto 0);
    signal conv53_469 : std_logic_vector(31 downto 0);
    signal conv56_482 : std_logic_vector(31 downto 0);
    signal conv61_491 : std_logic_vector(31 downto 0);
    signal conv63_495 : std_logic_vector(31 downto 0);
    signal conv65_499 : std_logic_vector(31 downto 0);
    signal conv71_513 : std_logic_vector(31 downto 0);
    signal conv74_517 : std_logic_vector(31 downto 0);
    signal conv82_539 : std_logic_vector(15 downto 0);
    signal conv85_552 : std_logic_vector(15 downto 0);
    signal conv8_344 : std_logic_vector(15 downto 0);
    signal conv91_564 : std_logic_vector(15 downto 0);
    signal conv94_577 : std_logic_vector(15 downto 0);
    signal exitcond23_1109 : std_logic_vector(0 downto 0);
    signal exitcond32_893 : std_logic_vector(0 downto 0);
    signal exitcond8_1556 : std_logic_vector(0 downto 0);
    signal exitcond_1229 : std_logic_vector(0 downto 0);
    signal inc234_1104 : std_logic_vector(31 downto 0);
    signal inc256_1224 : std_logic_vector(31 downto 0);
    signal inc416_1551 : std_logic_vector(31 downto 0);
    signal inc_888 : std_logic_vector(31 downto 0);
    signal ix_x0431_729 : std_logic_vector(31 downto 0);
    signal ix_x1427_945 : std_logic_vector(31 downto 0);
    signal ix_x2423_1197 : std_logic_vector(31 downto 0);
    signal ix_x3420_1427 : std_logic_vector(31 downto 0);
    signal mul241_1135 : std_logic_vector(31 downto 0);
    signal mul244_1140 : std_logic_vector(31 downto 0);
    signal mul66_509 : std_logic_vector(31 downto 0);
    signal mul72_522 : std_logic_vector(31 downto 0);
    signal mul75_527 : std_logic_vector(31 downto 0);
    signal mul78_532 : std_logic_vector(31 downto 0);
    signal mul_504 : std_logic_vector(31 downto 0);
    signal ptr_deref_1096_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1096_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1096_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1096_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1096_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1096_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1215_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1215_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1215_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1215_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1215_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1215_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1446_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1446_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1446_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1446_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1446_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_880_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_880_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_880_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_880_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_880_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_880_word_offset_0 : std_logic_vector(15 downto 0);
    signal shl101_595 : std_logic_vector(15 downto 0);
    signal shl110_620 : std_logic_vector(15 downto 0);
    signal shl119_645 : std_logic_vector(15 downto 0);
    signal shl132_758 : std_logic_vector(63 downto 0);
    signal shl138_776 : std_logic_vector(63 downto 0);
    signal shl144_794 : std_logic_vector(63 downto 0);
    signal shl150_812 : std_logic_vector(63 downto 0);
    signal shl156_830 : std_logic_vector(63 downto 0);
    signal shl162_848 : std_logic_vector(63 downto 0);
    signal shl168_866 : std_logic_vector(63 downto 0);
    signal shl188_974 : std_logic_vector(63 downto 0);
    signal shl18_375 : std_logic_vector(15 downto 0);
    signal shl194_992 : std_logic_vector(63 downto 0);
    signal shl200_1010 : std_logic_vector(63 downto 0);
    signal shl206_1028 : std_logic_vector(63 downto 0);
    signal shl212_1046 : std_logic_vector(63 downto 0);
    signal shl218_1064 : std_logic_vector(63 downto 0);
    signal shl224_1082 : std_logic_vector(63 downto 0);
    signal shl27_400 : std_logic_vector(31 downto 0);
    signal shl36_425 : std_logic_vector(15 downto 0);
    signal shl45_450 : std_logic_vector(15 downto 0);
    signal shl54_475 : std_logic_vector(31 downto 0);
    signal shl83_545 : std_logic_vector(15 downto 0);
    signal shl92_570 : std_logic_vector(15 downto 0);
    signal shl9_350 : std_logic_vector(15 downto 0);
    signal shl_325 : std_logic_vector(15 downto 0);
    signal shr282_1287 : std_logic_vector(63 downto 0);
    signal shr288_1297 : std_logic_vector(63 downto 0);
    signal shr294_1307 : std_logic_vector(63 downto 0);
    signal shr300_1317 : std_logic_vector(63 downto 0);
    signal shr306_1327 : std_logic_vector(63 downto 0);
    signal shr312_1337 : std_logic_vector(63 downto 0);
    signal shr318_1347 : std_logic_vector(63 downto 0);
    signal shr357_1457 : std_logic_vector(63 downto 0);
    signal shr363_1467 : std_logic_vector(63 downto 0);
    signal shr369_1477 : std_logic_vector(63 downto 0);
    signal shr375_1487 : std_logic_vector(63 downto 0);
    signal shr381_1497 : std_logic_vector(63 downto 0);
    signal shr387_1507 : std_logic_vector(63 downto 0);
    signal shr393_1517 : std_logic_vector(63 downto 0);
    signal sub_1276 : std_logic_vector(63 downto 0);
    signal tmp10_1161 : std_logic_vector(31 downto 0);
    signal tmp11_1166 : std_logic_vector(31 downto 0);
    signal tmp12_1170 : std_logic_vector(31 downto 0);
    signal tmp13_1175 : std_logic_vector(31 downto 0);
    signal tmp14_1181 : std_logic_vector(31 downto 0);
    signal tmp15_1187 : std_logic_vector(0 downto 0);
    signal tmp16_909 : std_logic_vector(31 downto 0);
    signal tmp17_914 : std_logic_vector(31 downto 0);
    signal tmp18_918 : std_logic_vector(31 downto 0);
    signal tmp19_923 : std_logic_vector(31 downto 0);
    signal tmp1_1391 : std_logic_vector(31 downto 0);
    signal tmp20_929 : std_logic_vector(31 downto 0);
    signal tmp21_935 : std_logic_vector(0 downto 0);
    signal tmp24_689 : std_logic_vector(31 downto 0);
    signal tmp25_693 : std_logic_vector(31 downto 0);
    signal tmp26_698 : std_logic_vector(31 downto 0);
    signal tmp27_702 : std_logic_vector(31 downto 0);
    signal tmp28_707 : std_logic_vector(31 downto 0);
    signal tmp29_713 : std_logic_vector(31 downto 0);
    signal tmp2_1396 : std_logic_vector(31 downto 0);
    signal tmp30_719 : std_logic_vector(0 downto 0);
    signal tmp350_1447 : std_logic_vector(63 downto 0);
    signal tmp3_1400 : std_logic_vector(31 downto 0);
    signal tmp448_905 : std_logic_vector(31 downto 0);
    signal tmp4_1405 : std_logic_vector(31 downto 0);
    signal tmp5_1411 : std_logic_vector(31 downto 0);
    signal tmp6_1417 : std_logic_vector(0 downto 0);
    signal tmp9_1157 : std_logic_vector(31 downto 0);
    signal tmp_1387 : std_logic_vector(31 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1026_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1044_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1062_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1102_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1179_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1192_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1201_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1203_wire : std_logic_vector(31 downto 0);
    signal type_cast_1217_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1222_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1245_wire : std_logic_vector(63 downto 0);
    signal type_cast_1260_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1262_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1269_wire : std_logic_vector(63 downto 0);
    signal type_cast_1285_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1295_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1305_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1315_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1325_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1335_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1345_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1409_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1415_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1422_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1431_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1433_wire : std_logic_vector(31 downto 0);
    signal type_cast_1455_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1465_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1475_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1485_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1495_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1505_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1515_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1549_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_323_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_348_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_373_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_398_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_423_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_473_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_543_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_568_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_593_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_618_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_643_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_661_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_711_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_717_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_733_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_735_wire : std_logic_vector(31 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_792_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_810_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_828_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_846_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_864_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_927_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_933_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_940_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_948_wire : std_logic_vector(31 downto 0);
    signal type_cast_951_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_972_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_990_wire_constant : std_logic_vector(63 downto 0);
    signal umax22_942 : std_logic_vector(31 downto 0);
    signal umax31_726 : std_logic_vector(31 downto 0);
    signal umax7_1424 : std_logic_vector(31 downto 0);
    signal umax_1194 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1211_constant_part_of_offset <= "1000000000000000";
    array_obj_ref_1211_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_1211_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_1211_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_1211_resized_base_address <= "0000000000000000";
    array_obj_ref_1441_constant_part_of_offset <= "1000000000000000";
    array_obj_ref_1441_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_1441_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_1441_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_1441_resized_base_address <= "0000000000000000";
    array_obj_ref_743_constant_part_of_offset <= "0000000000000000";
    array_obj_ref_743_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_743_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_743_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_743_resized_base_address <= "0000000000000000";
    array_obj_ref_959_constant_part_of_offset <= "0100000000000000";
    array_obj_ref_959_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_959_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_959_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_959_resized_base_address <= "0000000000000000";
    ptr_deref_1096_word_offset_0 <= "0000000000000000";
    ptr_deref_1215_word_offset_0 <= "0000000000000000";
    ptr_deref_1446_word_offset_0 <= "0000000000000000";
    ptr_deref_880_word_offset_0 <= "0000000000000000";
    type_cast_1008_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1026_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1044_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1062_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1080_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1102_wire_constant <= "00000000000000000000000000000001";
    type_cast_1144_wire_constant <= "00000000000000000000000000000111";
    type_cast_1179_wire_constant <= "00000000000000000000000000000011";
    type_cast_1185_wire_constant <= "00000000000000000000000000000001";
    type_cast_1192_wire_constant <= "00000000000000000000000000000001";
    type_cast_1201_wire_constant <= "00000000000000000000000000000000";
    type_cast_1217_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1222_wire_constant <= "00000000000000000000000000000001";
    type_cast_1260_wire_constant <= "00000000";
    type_cast_1262_wire_constant <= "00000010";
    type_cast_1285_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1295_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1305_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1315_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1325_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1335_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1345_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1409_wire_constant <= "00000000000000000000000000000011";
    type_cast_1415_wire_constant <= "00000000000000000000000000000001";
    type_cast_1422_wire_constant <= "00000000000000000000000000000001";
    type_cast_1431_wire_constant <= "00000000000000000000000000000000";
    type_cast_1455_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1465_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1475_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1485_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1495_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1505_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1515_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1549_wire_constant <= "00000000000000000000000000000001";
    type_cast_323_wire_constant <= "0000000000001000";
    type_cast_348_wire_constant <= "0000000000001000";
    type_cast_373_wire_constant <= "0000000000001000";
    type_cast_398_wire_constant <= "00000000000000000000000000001000";
    type_cast_423_wire_constant <= "0000000000001000";
    type_cast_448_wire_constant <= "0000000000001000";
    type_cast_473_wire_constant <= "00000000000000000000000000001000";
    type_cast_543_wire_constant <= "0000000000001000";
    type_cast_568_wire_constant <= "0000000000001000";
    type_cast_593_wire_constant <= "0000000000001000";
    type_cast_618_wire_constant <= "0000000000001000";
    type_cast_643_wire_constant <= "0000000000001000";
    type_cast_661_wire_constant <= "00000000000000000000000000000111";
    type_cast_676_wire_constant <= "00000000000000000000000000000111";
    type_cast_711_wire_constant <= "00000000000000000000000000000011";
    type_cast_717_wire_constant <= "00000000000000000000000000000001";
    type_cast_724_wire_constant <= "00000000000000000000000000000001";
    type_cast_733_wire_constant <= "00000000000000000000000000000000";
    type_cast_756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_774_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_792_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_810_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_828_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_846_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_864_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_886_wire_constant <= "00000000000000000000000000000001";
    type_cast_927_wire_constant <= "00000000000000000000000000000011";
    type_cast_933_wire_constant <= "00000000000000000000000000000001";
    type_cast_940_wire_constant <= "00000000000000000000000000000001";
    type_cast_951_wire_constant <= "00000000000000000000000000000000";
    type_cast_972_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_990_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    phi_stmt_1197: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1201_wire_constant & type_cast_1203_wire;
      req <= phi_stmt_1197_req_0 & phi_stmt_1197_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1197",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1197_ack_0,
          idata => idata,
          odata => ix_x2423_1197,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1197
    phi_stmt_1427: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1431_wire_constant & type_cast_1433_wire;
      req <= phi_stmt_1427_req_0 & phi_stmt_1427_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1427",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1427_ack_0,
          idata => idata,
          odata => ix_x3420_1427,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1427
    phi_stmt_729: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_733_wire_constant & type_cast_735_wire;
      req <= phi_stmt_729_req_0 & phi_stmt_729_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_729",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_729_ack_0,
          idata => idata,
          odata => ix_x0431_729,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_729
    phi_stmt_945: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_948_wire & type_cast_951_wire_constant;
      req <= phi_stmt_945_req_0 & phi_stmt_945_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_945",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_945_ack_0,
          idata => idata,
          odata => ix_x1427_945,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_945
    -- flow-through select operator MUX_1193_inst
    umax_1194 <= tmp14_1181 when (tmp15_1187(0) /=  '0') else type_cast_1192_wire_constant;
    -- flow-through select operator MUX_1423_inst
    umax7_1424 <= tmp5_1411 when (tmp6_1417(0) /=  '0') else type_cast_1422_wire_constant;
    -- flow-through select operator MUX_725_inst
    umax31_726 <= tmp29_713 when (tmp30_719(0) /=  '0') else type_cast_724_wire_constant;
    -- flow-through select operator MUX_941_inst
    umax22_942 <= tmp20_929 when (tmp21_935(0) /=  '0') else type_cast_940_wire_constant;
    addr_of_1212_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1212_final_reg_req_0;
      addr_of_1212_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1212_final_reg_req_1;
      addr_of_1212_final_reg_ack_1<= rack(0);
      addr_of_1212_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1212_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1211_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx253_1213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1442_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1442_final_reg_req_0;
      addr_of_1442_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1442_final_reg_req_1;
      addr_of_1442_final_reg_ack_1<= rack(0);
      addr_of_1442_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1442_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1441_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx349_1443,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_744_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_744_final_reg_req_0;
      addr_of_744_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_744_final_reg_req_1;
      addr_of_744_final_reg_ack_1<= rack(0);
      addr_of_744_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_744_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_743_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_745,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_960_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_960_final_reg_req_0;
      addr_of_960_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_960_final_reg_req_1;
      addr_of_960_final_reg_ack_1<= rack(0);
      addr_of_960_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_960_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_959_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx231_961,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1016_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1016_inst_req_0;
      type_cast_1016_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1016_inst_req_1;
      type_cast_1016_inst_ack_1<= rack(0);
      type_cast_1016_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1016_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call201_1013,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv203_1017,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1034_inst_req_0;
      type_cast_1034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1034_inst_req_1;
      type_cast_1034_inst_ack_1<= rack(0);
      type_cast_1034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call207_1031,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv209_1035,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1052_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1052_inst_req_0;
      type_cast_1052_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1052_inst_req_1;
      type_cast_1052_inst_ack_1<= rack(0);
      type_cast_1052_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1052_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call213_1049,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv215_1053,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1070_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1070_inst_req_0;
      type_cast_1070_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1070_inst_req_1;
      type_cast_1070_inst_ack_1<= rack(0);
      type_cast_1070_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1070_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call219_1067,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv221_1071,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1088_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1088_inst_req_0;
      type_cast_1088_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1088_inst_req_1;
      type_cast_1088_inst_ack_1<= rack(0);
      type_cast_1088_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1088_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call225_1085,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv227_1089,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1121_inst_req_0;
      type_cast_1121_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1121_inst_req_1;
      type_cast_1121_inst_ack_1<= rack(0);
      type_cast_1121_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1121_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add104_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv238_1122,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1125_inst_req_0;
      type_cast_1125_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1125_inst_req_1;
      type_cast_1125_inst_ack_1<= rack(0);
      type_cast_1125_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1125_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add113_632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv240_1126,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1129_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1129_inst_req_0;
      type_cast_1129_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1129_inst_req_1;
      type_cast_1129_inst_ack_1<= rack(0);
      type_cast_1129_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1129_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add122_657,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv243_1130,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1156_inst_req_0;
      type_cast_1156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1156_inst_req_1;
      type_cast_1156_inst_ack_1<= rack(0);
      type_cast_1156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add113_632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp9_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1160_inst_req_0;
      type_cast_1160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1160_inst_req_1;
      type_cast_1160_inst_ack_1<= rack(0);
      type_cast_1160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add104_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10_1161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1169_inst_req_0;
      type_cast_1169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1169_inst_req_1;
      type_cast_1169_inst_ack_1<= rack(0);
      type_cast_1169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add122_657,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_1170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1203_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1203_inst_req_0;
      type_cast_1203_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1203_inst_req_1;
      type_cast_1203_inst_ack_1<= rack(0);
      type_cast_1203_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1203_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc256_1224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1203_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1246_inst_req_0;
      type_cast_1246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1246_inst_req_1;
      type_cast_1246_inst_ack_1<= rack(0);
      type_cast_1246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1246_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1245_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv260_1247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1270_inst_req_0;
      type_cast_1270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1270_inst_req_1;
      type_cast_1270_inst_ack_1<= rack(0);
      type_cast_1270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1269_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv273_1271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1280_inst_req_0;
      type_cast_1280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1280_inst_req_1;
      type_cast_1280_inst_ack_1<= rack(0);
      type_cast_1280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv279_1281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1290_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1290_inst_req_0;
      type_cast_1290_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1290_inst_req_1;
      type_cast_1290_inst_ack_1<= rack(0);
      type_cast_1290_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1290_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr282_1287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv285_1291,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1300_inst_req_0;
      type_cast_1300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1300_inst_req_1;
      type_cast_1300_inst_ack_1<= rack(0);
      type_cast_1300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1300_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr288_1297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv291_1301,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1310_inst_req_0;
      type_cast_1310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1310_inst_req_1;
      type_cast_1310_inst_ack_1<= rack(0);
      type_cast_1310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr294_1307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv297_1311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1320_inst_req_0;
      type_cast_1320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1320_inst_req_1;
      type_cast_1320_inst_ack_1<= rack(0);
      type_cast_1320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr300_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv303_1321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1330_inst_req_0;
      type_cast_1330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1330_inst_req_1;
      type_cast_1330_inst_ack_1<= rack(0);
      type_cast_1330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr306_1327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv309_1331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1340_inst_req_0;
      type_cast_1340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1340_inst_req_1;
      type_cast_1340_inst_ack_1<= rack(0);
      type_cast_1340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr312_1337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv315_1341,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1350_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1350_inst_req_0;
      type_cast_1350_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1350_inst_req_1;
      type_cast_1350_inst_ack_1<= rack(0);
      type_cast_1350_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1350_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr318_1347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv321_1351,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1386_inst_req_0;
      type_cast_1386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1386_inst_req_1;
      type_cast_1386_inst_ack_1<= rack(0);
      type_cast_1386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add113_632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_1387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1390_inst_req_0;
      type_cast_1390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1390_inst_req_1;
      type_cast_1390_inst_ack_1<= rack(0);
      type_cast_1390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add104_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_1391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1399_inst_req_0;
      type_cast_1399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1399_inst_req_1;
      type_cast_1399_inst_ack_1<= rack(0);
      type_cast_1399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1399_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add122_657,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1433_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1433_inst_req_0;
      type_cast_1433_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1433_inst_req_1;
      type_cast_1433_inst_ack_1<= rack(0);
      type_cast_1433_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1433_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc416_1551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1433_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1450_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1450_inst_req_0;
      type_cast_1450_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1450_inst_req_1;
      type_cast_1450_inst_ack_1<= rack(0);
      type_cast_1450_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1450_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp350_1447,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv354_1451,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1460_inst_req_0;
      type_cast_1460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1460_inst_req_1;
      type_cast_1460_inst_ack_1<= rack(0);
      type_cast_1460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr357_1457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv360_1461,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1470_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1470_inst_req_0;
      type_cast_1470_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1470_inst_req_1;
      type_cast_1470_inst_ack_1<= rack(0);
      type_cast_1470_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1470_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr363_1467,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv366_1471,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1480_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1480_inst_req_0;
      type_cast_1480_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1480_inst_req_1;
      type_cast_1480_inst_ack_1<= rack(0);
      type_cast_1480_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1480_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr369_1477,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv372_1481,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1490_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1490_inst_req_0;
      type_cast_1490_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1490_inst_req_1;
      type_cast_1490_inst_ack_1<= rack(0);
      type_cast_1490_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1490_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr375_1487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv378_1491,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1500_inst_req_0;
      type_cast_1500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1500_inst_req_1;
      type_cast_1500_inst_ack_1<= rack(0);
      type_cast_1500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr381_1497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv384_1501,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1510_inst_req_0;
      type_cast_1510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1510_inst_req_1;
      type_cast_1510_inst_ack_1<= rack(0);
      type_cast_1510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr387_1507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv390_1511,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1520_inst_req_0;
      type_cast_1520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1520_inst_req_1;
      type_cast_1520_inst_ack_1<= rack(0);
      type_cast_1520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr393_1517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv396_1521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_318_inst_req_0;
      type_cast_318_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_318_inst_req_1;
      type_cast_318_inst_ack_1<= rack(0);
      type_cast_318_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_318_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_319,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_331_inst_req_0;
      type_cast_331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_331_inst_req_1;
      type_cast_331_inst_ack_1<= rack(0);
      type_cast_331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_328,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_343_inst_req_0;
      type_cast_343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_343_inst_req_1;
      type_cast_343_inst_ack_1<= rack(0);
      type_cast_343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_344,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_356_inst_req_0;
      type_cast_356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_356_inst_req_1;
      type_cast_356_inst_ack_1<= rack(0);
      type_cast_356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_353,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_368_inst_req_0;
      type_cast_368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_368_inst_req_1;
      type_cast_368_inst_ack_1<= rack(0);
      type_cast_368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_381_inst_req_0;
      type_cast_381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_381_inst_req_1;
      type_cast_381_inst_ack_1<= rack(0);
      type_cast_381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_381_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_393_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_393_inst_req_0;
      type_cast_393_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_393_inst_req_1;
      type_cast_393_inst_ack_1<= rack(0);
      type_cast_393_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_393_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_394,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_406_inst_req_0;
      type_cast_406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_406_inst_req_1;
      type_cast_406_inst_ack_1<= rack(0);
      type_cast_406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_403,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_418_inst_req_0;
      type_cast_418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_418_inst_req_1;
      type_cast_418_inst_ack_1<= rack(0);
      type_cast_418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_431_inst_req_0;
      type_cast_431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_431_inst_req_1;
      type_cast_431_inst_ack_1<= rack(0);
      type_cast_431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_428,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_432,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_443_inst_req_0;
      type_cast_443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_443_inst_req_1;
      type_cast_443_inst_ack_1<= rack(0);
      type_cast_443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_456_inst_req_0;
      type_cast_456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_456_inst_req_1;
      type_cast_456_inst_ack_1<= rack(0);
      type_cast_456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_457,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_468_inst_req_0;
      type_cast_468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_468_inst_req_1;
      type_cast_468_inst_ack_1<= rack(0);
      type_cast_468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_468_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_465,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_469,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_481_inst_req_0;
      type_cast_481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_481_inst_req_1;
      type_cast_481_inst_ack_1<= rack(0);
      type_cast_481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_482,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_490_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_490_inst_req_0;
      type_cast_490_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_490_inst_req_1;
      type_cast_490_inst_ack_1<= rack(0);
      type_cast_490_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_490_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_491,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_494_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_494_inst_req_0;
      type_cast_494_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_494_inst_req_1;
      type_cast_494_inst_ack_1<= rack(0);
      type_cast_494_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_494_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_362,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_495,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_498_inst_req_0;
      type_cast_498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_498_inst_req_1;
      type_cast_498_inst_ack_1<= rack(0);
      type_cast_498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_512_inst_req_0;
      type_cast_512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_512_inst_req_1;
      type_cast_512_inst_ack_1<= rack(0);
      type_cast_512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_437,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_513,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_516_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_516_inst_req_0;
      type_cast_516_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_516_inst_req_1;
      type_cast_516_inst_ack_1<= rack(0);
      type_cast_516_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_516_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_517,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_538_inst_req_1;
      type_cast_538_inst_ack_1<= rack(0);
      type_cast_538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call79_535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_551_inst_req_0;
      type_cast_551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_551_inst_req_1;
      type_cast_551_inst_ack_1<= rack(0);
      type_cast_551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_563_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_563_inst_req_0;
      type_cast_563_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_563_inst_req_1;
      type_cast_563_inst_ack_1<= rack(0);
      type_cast_563_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_563_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_560,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_564,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_576_inst_req_0;
      type_cast_576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_576_inst_req_1;
      type_cast_576_inst_ack_1<= rack(0);
      type_cast_576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_573,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_588_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_588_inst_req_0;
      type_cast_588_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_588_inst_req_1;
      type_cast_588_inst_ack_1<= rack(0);
      type_cast_588_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_588_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_589,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_601_inst_req_0;
      type_cast_601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_601_inst_req_1;
      type_cast_601_inst_ack_1<= rack(0);
      type_cast_601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call102_598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_613_inst_req_0;
      type_cast_613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_613_inst_req_1;
      type_cast_613_inst_ack_1<= rack(0);
      type_cast_613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_626_inst_req_0;
      type_cast_626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_626_inst_req_1;
      type_cast_626_inst_ack_1<= rack(0);
      type_cast_626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_638_inst_req_0;
      type_cast_638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_638_inst_req_1;
      type_cast_638_inst_ack_1<= rack(0);
      type_cast_638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_638_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_635,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_639,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_651_inst_req_0;
      type_cast_651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_651_inst_req_1;
      type_cast_651_inst_ack_1<= rack(0);
      type_cast_651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_651_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call120_648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_652,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_688_inst_req_0;
      type_cast_688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_688_inst_req_1;
      type_cast_688_inst_ack_1<= rack(0);
      type_cast_688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_362,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_692_inst_req_0;
      type_cast_692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_692_inst_req_1;
      type_cast_692_inst_ack_1<= rack(0);
      type_cast_692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_692_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp25_693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_701_inst_req_0;
      type_cast_701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_701_inst_req_1;
      type_cast_701_inst_ack_1<= rack(0);
      type_cast_701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp27_702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_735_inst_req_0;
      type_cast_735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_735_inst_req_1;
      type_cast_735_inst_ack_1<= rack(0);
      type_cast_735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_888,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_735_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_751_inst_req_1;
      type_cast_751_inst_ack_1<= rack(0);
      type_cast_751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_764_inst_req_0;
      type_cast_764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_764_inst_req_1;
      type_cast_764_inst_ack_1<= rack(0);
      type_cast_764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_782_inst_req_0;
      type_cast_782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_782_inst_req_1;
      type_cast_782_inst_ack_1<= rack(0);
      type_cast_782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call139_779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_800_inst_req_0;
      type_cast_800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_800_inst_req_1;
      type_cast_800_inst_ack_1<= rack(0);
      type_cast_800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_818_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_818_inst_req_0;
      type_cast_818_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_818_inst_req_1;
      type_cast_818_inst_ack_1<= rack(0);
      type_cast_818_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_818_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call151_815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_819,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_836_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_836_inst_req_0;
      type_cast_836_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_836_inst_req_1;
      type_cast_836_inst_ack_1<= rack(0);
      type_cast_836_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_836_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_837,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack(0);
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_851,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_872_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_872_inst_req_0;
      type_cast_872_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_872_inst_req_1;
      type_cast_872_inst_ack_1<= rack(0);
      type_cast_872_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_872_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_869,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_873,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_908_inst_req_0;
      type_cast_908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_908_inst_req_1;
      type_cast_908_inst_ack_1<= rack(0);
      type_cast_908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_908_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_437,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_909,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_917_inst_req_0;
      type_cast_917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_917_inst_req_1;
      type_cast_917_inst_ack_1<= rack(0);
      type_cast_917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp18_918,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_948_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_948_inst_req_0;
      type_cast_948_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_948_inst_req_1;
      type_cast_948_inst_ack_1<= rack(0);
      type_cast_948_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_948_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc234_1104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_948_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_967_inst_req_0;
      type_cast_967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_967_inst_req_1;
      type_cast_967_inst_ack_1<= rack(0);
      type_cast_967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call185_964,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv186_968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_980_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_980_inst_req_0;
      type_cast_980_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_980_inst_req_1;
      type_cast_980_inst_ack_1<= rack(0);
      type_cast_980_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_980_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call189_977,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_981,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_998_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_998_inst_req_0;
      type_cast_998_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_998_inst_req_1;
      type_cast_998_inst_ack_1<= rack(0);
      type_cast_998_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_998_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call195_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv197_999,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1211_index_2_rename
    process(R_ix_x2423_1210_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x2423_1210_resized;
      ov(15 downto 0) := iv;
      R_ix_x2423_1210_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1211_index_2_resize
    process(ix_x2423_1197) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x2423_1197;
      ov := iv(15 downto 0);
      R_ix_x2423_1210_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1211_root_address_inst
    process(array_obj_ref_1211_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1211_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_1211_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_index_2_rename
    process(R_ix_x3420_1440_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x3420_1440_resized;
      ov(15 downto 0) := iv;
      R_ix_x3420_1440_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_index_2_resize
    process(ix_x3420_1427) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x3420_1427;
      ov := iv(15 downto 0);
      R_ix_x3420_1440_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_root_address_inst
    process(array_obj_ref_1441_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1441_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_1441_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_743_index_2_rename
    process(R_ix_x0431_742_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0431_742_resized;
      ov(15 downto 0) := iv;
      R_ix_x0431_742_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_743_index_2_resize
    process(ix_x0431_729) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0431_729;
      ov := iv(15 downto 0);
      R_ix_x0431_742_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_743_root_address_inst
    process(array_obj_ref_743_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_743_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_743_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_959_index_2_rename
    process(R_ix_x1427_958_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1427_958_resized;
      ov(15 downto 0) := iv;
      R_ix_x1427_958_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_959_index_2_resize
    process(ix_x1427_945) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1427_945;
      ov := iv(15 downto 0);
      R_ix_x1427_958_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_959_root_address_inst
    process(array_obj_ref_959_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_959_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_959_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_addr_0
    process(ptr_deref_1096_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1096_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_1096_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_base_resize
    process(arrayidx231_961) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx231_961;
      ov := iv(15 downto 0);
      ptr_deref_1096_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_gather_scatter
    process(add228_1094) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add228_1094;
      ov(63 downto 0) := iv;
      ptr_deref_1096_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_root_address_inst
    process(ptr_deref_1096_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1096_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_1096_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1215_addr_0
    process(ptr_deref_1215_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1215_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_1215_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1215_base_resize
    process(arrayidx253_1213) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx253_1213;
      ov := iv(15 downto 0);
      ptr_deref_1215_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1215_gather_scatter
    process(type_cast_1217_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1217_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1215_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1215_root_address_inst
    process(ptr_deref_1215_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1215_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_1215_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1446_addr_0
    process(ptr_deref_1446_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1446_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_1446_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1446_base_resize
    process(arrayidx349_1443) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx349_1443;
      ov := iv(15 downto 0);
      ptr_deref_1446_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1446_gather_scatter
    process(ptr_deref_1446_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1446_data_0;
      ov(63 downto 0) := iv;
      tmp350_1447 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1446_root_address_inst
    process(ptr_deref_1446_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1446_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_1446_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_addr_0
    process(ptr_deref_880_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_880_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_880_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_base_resize
    process(arrayidx_745) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_745;
      ov := iv(15 downto 0);
      ptr_deref_880_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_gather_scatter
    process(add172_878) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add172_878;
      ov(63 downto 0) := iv;
      ptr_deref_880_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_root_address_inst
    process(ptr_deref_880_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_880_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_880_root_address <= ov(15 downto 0);
      --
    end process;
    if_stmt_1110_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond23_1109;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1110_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1110_branch_req_0,
          ack0 => if_stmt_1110_branch_ack_0,
          ack1 => if_stmt_1110_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1147_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp249422_1146;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1147_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1147_branch_req_0,
          ack0 => if_stmt_1147_branch_ack_0,
          ack1 => if_stmt_1147_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1230_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1229;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1230_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1230_branch_req_0,
          ack0 => if_stmt_1230_branch_ack_0,
          ack1 => if_stmt_1230_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1377_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp249422_1146;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1377_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1377_branch_req_0,
          ack0 => if_stmt_1377_branch_ack_0,
          ack1 => if_stmt_1377_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1557_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond8_1556;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1557_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1557_branch_req_0,
          ack0 => if_stmt_1557_branch_ack_0,
          ack1 => if_stmt_1557_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_664_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp430_663;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_664_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_664_branch_req_0,
          ack0 => if_stmt_664_branch_ack_0,
          ack1 => if_stmt_664_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_679_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp180426_678;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_679_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_679_branch_req_0,
          ack0 => if_stmt_679_branch_ack_0,
          ack1 => if_stmt_679_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_894_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond32_893;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_894_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_894_branch_req_0,
          ack0 => if_stmt_894_branch_ack_0,
          ack1 => if_stmt_894_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1103_inst
    process(ix_x1427_945) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x1427_945, type_cast_1102_wire_constant, tmp_var);
      inc234_1104 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1223_inst
    process(ix_x2423_1197) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x2423_1197, type_cast_1222_wire_constant, tmp_var);
      inc256_1224 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1550_inst
    process(ix_x3420_1427) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x3420_1427, type_cast_1549_wire_constant, tmp_var);
      inc416_1551 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_887_inst
    process(ix_x0431_729) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x0431_729, type_cast_886_wire_constant, tmp_var);
      inc_888 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1108_inst
    process(inc234_1104, umax22_942) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc234_1104, umax22_942, tmp_var);
      exitcond23_1109 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1228_inst
    process(inc256_1224, umax_1194) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc256_1224, umax_1194, tmp_var);
      exitcond_1229 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1555_inst
    process(inc416_1551, umax7_1424) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc416_1551, umax7_1424, tmp_var);
      exitcond8_1556 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_892_inst
    process(inc_888, umax31_726) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_888, umax31_726, tmp_var);
      exitcond32_893 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1180_inst
    process(tmp13_1175) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp13_1175, type_cast_1179_wire_constant, tmp_var);
      tmp14_1181 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1410_inst
    process(tmp4_1405) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1405, type_cast_1409_wire_constant, tmp_var);
      tmp5_1411 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_712_inst
    process(tmp28_707) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp28_707, type_cast_711_wire_constant, tmp_var);
      tmp29_713 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_928_inst
    process(tmp19_923) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp19_923, type_cast_927_wire_constant, tmp_var);
      tmp20_929 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1286_inst
    process(sub_1276) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1276, type_cast_1285_wire_constant, tmp_var);
      shr282_1287 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1296_inst
    process(sub_1276) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1276, type_cast_1295_wire_constant, tmp_var);
      shr288_1297 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1306_inst
    process(sub_1276) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1276, type_cast_1305_wire_constant, tmp_var);
      shr294_1307 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1316_inst
    process(sub_1276) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1276, type_cast_1315_wire_constant, tmp_var);
      shr300_1317 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1326_inst
    process(sub_1276) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1276, type_cast_1325_wire_constant, tmp_var);
      shr306_1327 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1336_inst
    process(sub_1276) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1276, type_cast_1335_wire_constant, tmp_var);
      shr312_1337 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1346_inst
    process(sub_1276) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1276, type_cast_1345_wire_constant, tmp_var);
      shr318_1347 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1456_inst
    process(tmp350_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp350_1447, type_cast_1455_wire_constant, tmp_var);
      shr357_1457 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1466_inst
    process(tmp350_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp350_1447, type_cast_1465_wire_constant, tmp_var);
      shr363_1467 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1476_inst
    process(tmp350_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp350_1447, type_cast_1475_wire_constant, tmp_var);
      shr369_1477 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1486_inst
    process(tmp350_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp350_1447, type_cast_1485_wire_constant, tmp_var);
      shr375_1487 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1496_inst
    process(tmp350_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp350_1447, type_cast_1495_wire_constant, tmp_var);
      shr381_1497 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1506_inst
    process(tmp350_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp350_1447, type_cast_1505_wire_constant, tmp_var);
      shr387_1507 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1516_inst
    process(tmp350_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp350_1447, type_cast_1515_wire_constant, tmp_var);
      shr393_1517 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1134_inst
    process(conv240_1126, conv238_1122) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv240_1126, conv238_1122, tmp_var);
      mul241_1135 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1139_inst
    process(mul241_1135, conv243_1130) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul241_1135, conv243_1130, tmp_var);
      mul244_1140 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1165_inst
    process(tmp9_1157, tmp10_1161) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1157, tmp10_1161, tmp_var);
      tmp11_1166 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1174_inst
    process(tmp11_1166, tmp12_1170) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_1166, tmp12_1170, tmp_var);
      tmp13_1175 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1395_inst
    process(tmp_1387, tmp1_1391) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1387, tmp1_1391, tmp_var);
      tmp2_1396 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1404_inst
    process(tmp2_1396, tmp3_1400) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_1396, tmp3_1400, tmp_var);
      tmp4_1405 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_503_inst
    process(conv63_495, conv61_491) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_495, conv61_491, tmp_var);
      mul_504 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_508_inst
    process(mul_504, conv65_499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_504, conv65_499, tmp_var);
      mul66_509 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_521_inst
    process(conv71_513, add30_412) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_513, add30_412, tmp_var);
      mul72_522 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_526_inst
    process(mul72_522, conv74_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul72_522, conv74_517, tmp_var);
      mul75_527 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_531_inst
    process(mul75_527, add57_487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul75_527, add57_487, tmp_var);
      mul78_532 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_697_inst
    process(tmp24_689, tmp25_693) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp24_689, tmp25_693, tmp_var);
      tmp26_698 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_706_inst
    process(tmp26_698, tmp27_702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp26_698, tmp27_702, tmp_var);
      tmp28_707 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_904_inst
    process(add30_412, add57_487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add30_412, add57_487, tmp_var);
      tmp448_905 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_913_inst
    process(tmp448_905, tmp16_909) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp448_905, tmp16_909, tmp_var);
      tmp17_914 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_922_inst
    process(tmp17_914, tmp18_918) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp17_914, tmp18_918, tmp_var);
      tmp19_923 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_336_inst
    process(shl_325, conv3_332) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_325, conv3_332, tmp_var);
      add_337 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_361_inst
    process(shl9_350, conv11_357) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_350, conv11_357, tmp_var);
      add12_362 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_386_inst
    process(shl18_375, conv20_382) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_375, conv20_382, tmp_var);
      add21_387 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_436_inst
    process(shl36_425, conv38_432) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_425, conv38_432, tmp_var);
      add39_437 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_461_inst
    process(shl45_450, conv47_457) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_450, conv47_457, tmp_var);
      add48_462 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_556_inst
    process(shl83_545, conv85_552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_545, conv85_552, tmp_var);
      add86_557 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_581_inst
    process(shl92_570, conv94_577) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_570, conv94_577, tmp_var);
      add95_582 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_606_inst
    process(shl101_595, conv103_602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl101_595, conv103_602, tmp_var);
      add104_607 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_631_inst
    process(shl110_620, conv112_627) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_620, conv112_627, tmp_var);
      add113_632 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_656_inst
    process(shl119_645, conv121_652) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl119_645, conv121_652, tmp_var);
      add122_657 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_411_inst
    process(shl27_400, conv29_407) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_400, conv29_407, tmp_var);
      add30_412 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_486_inst
    process(shl54_475, conv56_482) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_475, conv56_482, tmp_var);
      add57_487 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1003_inst
    process(shl194_992, conv197_999) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl194_992, conv197_999, tmp_var);
      add198_1004 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1021_inst
    process(shl200_1010, conv203_1017) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl200_1010, conv203_1017, tmp_var);
      add204_1022 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1039_inst
    process(shl206_1028, conv209_1035) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl206_1028, conv209_1035, tmp_var);
      add210_1040 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1057_inst
    process(shl212_1046, conv215_1053) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl212_1046, conv215_1053, tmp_var);
      add216_1058 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1075_inst
    process(shl218_1064, conv221_1071) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl218_1064, conv221_1071, tmp_var);
      add222_1076 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1093_inst
    process(shl224_1082, conv227_1089) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl224_1082, conv227_1089, tmp_var);
      add228_1094 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_769_inst
    process(shl132_758, conv135_765) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_758, conv135_765, tmp_var);
      add136_770 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_787_inst
    process(shl138_776, conv141_783) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl138_776, conv141_783, tmp_var);
      add142_788 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_805_inst
    process(shl144_794, conv147_801) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_794, conv147_801, tmp_var);
      add148_806 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_823_inst
    process(shl150_812, conv153_819) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl150_812, conv153_819, tmp_var);
      add154_824 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_841_inst
    process(shl156_830, conv159_837) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_830, conv159_837, tmp_var);
      add160_842 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_859_inst
    process(shl162_848, conv165_855) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_848, conv165_855, tmp_var);
      add166_860 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_877_inst
    process(shl168_866, conv171_873) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_866, conv171_873, tmp_var);
      add172_878 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_985_inst
    process(shl188_974, conv191_981) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl188_974, conv191_981, tmp_var);
      add192_986 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_324_inst
    process(conv1_319) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_319, type_cast_323_wire_constant, tmp_var);
      shl_325 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_349_inst
    process(conv8_344) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_344, type_cast_348_wire_constant, tmp_var);
      shl9_350 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_374_inst
    process(conv17_369) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_369, type_cast_373_wire_constant, tmp_var);
      shl18_375 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_424_inst
    process(conv35_419) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_419, type_cast_423_wire_constant, tmp_var);
      shl36_425 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_449_inst
    process(conv44_444) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_444, type_cast_448_wire_constant, tmp_var);
      shl45_450 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_544_inst
    process(conv82_539) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv82_539, type_cast_543_wire_constant, tmp_var);
      shl83_545 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_569_inst
    process(conv91_564) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_564, type_cast_568_wire_constant, tmp_var);
      shl92_570 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_594_inst
    process(conv100_589) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv100_589, type_cast_593_wire_constant, tmp_var);
      shl101_595 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_619_inst
    process(conv109_614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv109_614, type_cast_618_wire_constant, tmp_var);
      shl110_620 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_644_inst
    process(conv118_639) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv118_639, type_cast_643_wire_constant, tmp_var);
      shl119_645 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_399_inst
    process(conv26_394) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_394, type_cast_398_wire_constant, tmp_var);
      shl27_400 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_474_inst
    process(conv53_469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_469, type_cast_473_wire_constant, tmp_var);
      shl54_475 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1009_inst
    process(add198_1004) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add198_1004, type_cast_1008_wire_constant, tmp_var);
      shl200_1010 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1027_inst
    process(add204_1022) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add204_1022, type_cast_1026_wire_constant, tmp_var);
      shl206_1028 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1045_inst
    process(add210_1040) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add210_1040, type_cast_1044_wire_constant, tmp_var);
      shl212_1046 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1063_inst
    process(add216_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add216_1058, type_cast_1062_wire_constant, tmp_var);
      shl218_1064 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1081_inst
    process(add222_1076) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add222_1076, type_cast_1080_wire_constant, tmp_var);
      shl224_1082 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_757_inst
    process(conv130_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv130_752, type_cast_756_wire_constant, tmp_var);
      shl132_758 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_775_inst
    process(add136_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add136_770, type_cast_774_wire_constant, tmp_var);
      shl138_776 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_793_inst
    process(add142_788) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add142_788, type_cast_792_wire_constant, tmp_var);
      shl144_794 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_811_inst
    process(add148_806) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add148_806, type_cast_810_wire_constant, tmp_var);
      shl150_812 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_829_inst
    process(add154_824) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add154_824, type_cast_828_wire_constant, tmp_var);
      shl156_830 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_847_inst
    process(add160_842) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_842, type_cast_846_wire_constant, tmp_var);
      shl162_848 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_865_inst
    process(add166_860) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_860, type_cast_864_wire_constant, tmp_var);
      shl168_866 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_973_inst
    process(conv186_968) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv186_968, type_cast_972_wire_constant, tmp_var);
      shl188_974 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_991_inst
    process(add192_986) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add192_986, type_cast_990_wire_constant, tmp_var);
      shl194_992 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1275_inst
    process(conv273_1271, conv260_1247) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv273_1271, conv260_1247, tmp_var);
      sub_1276 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1145_inst
    process(mul244_1140) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul244_1140, type_cast_1144_wire_constant, tmp_var);
      cmp249422_1146 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1186_inst
    process(tmp14_1181) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp14_1181, type_cast_1185_wire_constant, tmp_var);
      tmp15_1187 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1416_inst
    process(tmp5_1411) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp5_1411, type_cast_1415_wire_constant, tmp_var);
      tmp6_1417 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_662_inst
    process(mul66_509) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_509, type_cast_661_wire_constant, tmp_var);
      cmp430_663 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_677_inst
    process(mul78_532) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul78_532, type_cast_676_wire_constant, tmp_var);
      cmp180426_678 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_718_inst
    process(tmp29_713) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp29_713, type_cast_717_wire_constant, tmp_var);
      tmp30_719 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_934_inst
    process(tmp20_929) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp20_929, type_cast_933_wire_constant, tmp_var);
      tmp21_935 <= tmp_var; --
    end process;
    -- shared split operator group (102) : array_obj_ref_1211_index_offset 
    ApIntAdd_group_102: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x2423_1210_scaled;
      array_obj_ref_1211_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1211_index_offset_req_0;
      array_obj_ref_1211_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1211_index_offset_req_1;
      array_obj_ref_1211_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_102_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_102_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_102",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : array_obj_ref_1441_index_offset 
    ApIntAdd_group_103: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x3420_1440_scaled;
      array_obj_ref_1441_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1441_index_offset_req_0;
      array_obj_ref_1441_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1441_index_offset_req_1;
      array_obj_ref_1441_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_103_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_103_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_103",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : array_obj_ref_743_index_offset 
    ApIntAdd_group_104: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0431_742_scaled;
      array_obj_ref_743_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_743_index_offset_req_0;
      array_obj_ref_743_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_743_index_offset_req_1;
      array_obj_ref_743_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_104_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_104_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_104",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- shared split operator group (105) : array_obj_ref_959_index_offset 
    ApIntAdd_group_105: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1427_958_scaled;
      array_obj_ref_959_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_959_index_offset_req_0;
      array_obj_ref_959_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_959_index_offset_req_1;
      array_obj_ref_959_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_105_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_105_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_105",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0100000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 105
    -- unary operator type_cast_1245_inst
    process(call259_1241) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call259_1241, tmp_var);
      type_cast_1245_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1269_inst
    process(call272_1266) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call272_1266, tmp_var);
      type_cast_1269_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1446_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1446_load_0_req_0;
      ptr_deref_1446_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1446_load_0_req_1;
      ptr_deref_1446_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1446_word_address_0;
      ptr_deref_1446_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(15 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1215_store_0 ptr_deref_1096_store_0 ptr_deref_880_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(47 downto 0);
      signal data_in: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1215_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1096_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_880_store_0_req_0;
      ptr_deref_1215_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1096_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_880_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1215_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1096_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_880_store_0_req_1;
      ptr_deref_1215_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1096_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_880_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1215_word_address_0 & ptr_deref_1096_word_address_0 & ptr_deref_880_word_address_0;
      data_in <= ptr_deref_1215_data_0 & ptr_deref_1096_data_0 & ptr_deref_880_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 16,
        data_width => 64,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(15 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_1012_inst RPIPE_ConvTranspose_input_pipe_414_inst RPIPE_ConvTranspose_input_pipe_402_inst RPIPE_ConvTranspose_input_pipe_364_inst RPIPE_ConvTranspose_input_pipe_389_inst RPIPE_ConvTranspose_input_pipe_427_inst RPIPE_ConvTranspose_input_pipe_1066_inst RPIPE_ConvTranspose_input_pipe_314_inst RPIPE_ConvTranspose_input_pipe_352_inst RPIPE_ConvTranspose_input_pipe_439_inst RPIPE_ConvTranspose_input_pipe_377_inst RPIPE_ConvTranspose_input_pipe_327_inst RPIPE_ConvTranspose_input_pipe_1030_inst RPIPE_ConvTranspose_input_pipe_452_inst RPIPE_ConvTranspose_input_pipe_1048_inst RPIPE_ConvTranspose_input_pipe_994_inst RPIPE_ConvTranspose_input_pipe_339_inst RPIPE_ConvTranspose_input_pipe_1084_inst RPIPE_ConvTranspose_input_pipe_547_inst RPIPE_ConvTranspose_input_pipe_534_inst RPIPE_ConvTranspose_input_pipe_584_inst RPIPE_ConvTranspose_input_pipe_477_inst RPIPE_ConvTranspose_input_pipe_464_inst RPIPE_ConvTranspose_input_pipe_572_inst RPIPE_ConvTranspose_input_pipe_976_inst RPIPE_ConvTranspose_input_pipe_559_inst RPIPE_ConvTranspose_input_pipe_963_inst RPIPE_ConvTranspose_input_pipe_597_inst RPIPE_ConvTranspose_input_pipe_609_inst RPIPE_ConvTranspose_input_pipe_622_inst RPIPE_ConvTranspose_input_pipe_634_inst RPIPE_ConvTranspose_input_pipe_647_inst RPIPE_ConvTranspose_input_pipe_747_inst RPIPE_ConvTranspose_input_pipe_760_inst RPIPE_ConvTranspose_input_pipe_778_inst RPIPE_ConvTranspose_input_pipe_796_inst RPIPE_ConvTranspose_input_pipe_814_inst RPIPE_ConvTranspose_input_pipe_832_inst RPIPE_ConvTranspose_input_pipe_850_inst RPIPE_ConvTranspose_input_pipe_868_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_1012_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_414_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_402_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_364_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_389_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_427_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_1066_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_314_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_352_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_439_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_377_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_327_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_1030_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_452_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_1048_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_994_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_339_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_1084_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_547_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_584_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_477_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_464_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_572_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_976_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_559_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_963_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_597_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_609_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_622_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_634_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_647_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_747_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_814_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_832_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_850_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_868_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_1012_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_414_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_402_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_364_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_389_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_427_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_1066_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_314_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_352_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_439_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_377_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_327_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_1030_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_452_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_1048_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_994_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_339_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_1084_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_547_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_584_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_477_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_464_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_572_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_976_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_559_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_963_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_597_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_609_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_622_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_634_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_647_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_747_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_814_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_832_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_850_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_868_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_1012_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_414_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_402_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_364_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_389_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_427_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_1066_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_314_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_352_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_439_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_377_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_327_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_1030_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_452_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_1048_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_994_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_339_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_1084_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_547_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_584_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_477_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_464_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_572_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_976_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_559_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_963_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_597_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_609_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_622_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_634_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_647_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_747_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_814_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_832_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_850_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_868_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_1012_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_414_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_402_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_364_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_389_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_427_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_1066_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_314_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_352_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_439_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_377_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_327_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_1030_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_452_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_1048_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_994_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_339_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_1084_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_547_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_584_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_477_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_464_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_572_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_976_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_559_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_963_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_597_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_609_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_622_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_634_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_647_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_747_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_814_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_832_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_850_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_868_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call201_1013 <= data_out(319 downto 312);
      call32_415 <= data_out(311 downto 304);
      call28_403 <= data_out(303 downto 296);
      call14_365 <= data_out(295 downto 288);
      call23_390 <= data_out(287 downto 280);
      call37_428 <= data_out(279 downto 272);
      call219_1067 <= data_out(271 downto 264);
      call_315 <= data_out(263 downto 256);
      call10_353 <= data_out(255 downto 248);
      call41_440 <= data_out(247 downto 240);
      call19_378 <= data_out(239 downto 232);
      call2_328 <= data_out(231 downto 224);
      call207_1031 <= data_out(223 downto 216);
      call46_453 <= data_out(215 downto 208);
      call213_1049 <= data_out(207 downto 200);
      call195_995 <= data_out(199 downto 192);
      call5_340 <= data_out(191 downto 184);
      call225_1085 <= data_out(183 downto 176);
      call84_548 <= data_out(175 downto 168);
      call79_535 <= data_out(167 downto 160);
      call97_585 <= data_out(159 downto 152);
      call55_478 <= data_out(151 downto 144);
      call50_465 <= data_out(143 downto 136);
      call93_573 <= data_out(135 downto 128);
      call189_977 <= data_out(127 downto 120);
      call88_560 <= data_out(119 downto 112);
      call185_964 <= data_out(111 downto 104);
      call102_598 <= data_out(103 downto 96);
      call106_610 <= data_out(95 downto 88);
      call111_623 <= data_out(87 downto 80);
      call115_635 <= data_out(79 downto 72);
      call120_648 <= data_out(71 downto 64);
      call129_748 <= data_out(63 downto 56);
      call133_761 <= data_out(55 downto 48);
      call139_779 <= data_out(47 downto 40);
      call145_797 <= data_out(39 downto 32);
      call151_815 <= data_out(31 downto 24);
      call157_833 <= data_out(23 downto 16);
      call163_851 <= data_out(15 downto 8);
      call169_869 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1540_inst WPIPE_ConvTranspose_output_pipe_1525_inst WPIPE_ConvTranspose_output_pipe_1352_inst WPIPE_ConvTranspose_output_pipe_1355_inst WPIPE_ConvTranspose_output_pipe_1370_inst WPIPE_ConvTranspose_output_pipe_1358_inst WPIPE_ConvTranspose_output_pipe_1528_inst WPIPE_ConvTranspose_output_pipe_1361_inst WPIPE_ConvTranspose_output_pipe_1373_inst WPIPE_ConvTranspose_output_pipe_1364_inst WPIPE_ConvTranspose_output_pipe_1367_inst WPIPE_ConvTranspose_output_pipe_1531_inst WPIPE_ConvTranspose_output_pipe_1537_inst WPIPE_ConvTranspose_output_pipe_1522_inst WPIPE_ConvTranspose_output_pipe_1543_inst WPIPE_ConvTranspose_output_pipe_1534_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1540_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1525_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1352_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1355_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1370_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1358_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1528_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1361_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1373_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1364_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1367_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1531_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1537_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1522_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1543_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1534_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1540_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1525_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1352_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1355_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1370_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1358_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1528_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1361_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1373_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1364_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1367_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1531_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1537_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1522_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1543_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1534_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1540_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1525_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1352_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1355_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1370_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1358_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1528_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1361_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1373_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1364_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1367_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1531_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1537_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1522_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1543_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1534_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1540_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1525_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1352_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1355_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1370_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1358_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1528_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1361_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1373_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1364_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1367_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1531_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1537_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1522_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1543_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1534_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv360_1461 & conv390_1511 & conv321_1351 & conv315_1341 & conv285_1291 & conv309_1331 & conv384_1501 & conv303_1321 & conv279_1281 & conv297_1311 & conv291_1301 & conv378_1491 & conv366_1471 & conv396_1521 & conv354_1451 & conv372_1481;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1241_call call_stmt_1266_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1241_call_req_0;
      reqL_unguarded(0) <= call_stmt_1266_call_req_0;
      call_stmt_1241_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1266_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1241_call_req_1;
      reqR_unguarded(0) <= call_stmt_1266_call_req_1;
      call_stmt_1241_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1266_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call259_1241 <= data_out(127 downto 64);
      call272_1266 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1263_call 
    ct_core_call_group_1: Block -- 
      signal data_in: std_logic_vector(175 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1263_call_req_0;
      call_stmt_1263_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1263_call_req_1;
      call_stmt_1263_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      ct_core_call_group_1_gI: SplitGuardInterface generic map(name => "ct_core_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add_337 & add12_362 & add21_387 & add39_437 & add48_462 & add104_607 & add113_632 & add122_657 & add86_557 & add95_582 & type_cast_1260_wire_constant & type_cast_1262_wire_constant;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 176,
        owidth => 176,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ct_core_call_reqs(0),
          ackR => ct_core_call_acks(0),
          dataR => ct_core_call_data(175 downto 0),
          tagR => ct_core_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => ct_core_return_acks(0), -- cross-over
          ackL => ct_core_return_reqs(0), -- cross-over
          tagL => ct_core_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ct_core is -- 
  generic (tag_length : integer); 
  port ( -- 
    inp_d0 : in  std_logic_vector(15 downto 0);
    inp_d1 : in  std_logic_vector(15 downto 0);
    inp_d2 : in  std_logic_vector(15 downto 0);
    ker_d1 : in  std_logic_vector(15 downto 0);
    ker_d2 : in  std_logic_vector(15 downto 0);
    out_d0 : in  std_logic_vector(15 downto 0);
    out_d1 : in  std_logic_vector(15 downto 0);
    out_d2 : in  std_logic_vector(15 downto 0);
    stride : in  std_logic_vector(15 downto 0);
    padding : in  std_logic_vector(15 downto 0);
    index1 : in  std_logic_vector(7 downto 0);
    index3 : in  std_logic_vector(7 downto 0);
    readModule1_call_reqs : out  std_logic_vector(0 downto 0);
    readModule1_call_acks : in   std_logic_vector(0 downto 0);
    readModule1_call_data : out  std_logic_vector(39 downto 0);
    readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
    readModule1_return_reqs : out  std_logic_vector(0 downto 0);
    readModule1_return_acks : in   std_logic_vector(0 downto 0);
    readModule1_return_data : in   std_logic_vector(63 downto 0);
    readModule1_return_tag :  in   std_logic_vector(0 downto 0);
    writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_call_acks : in   std_logic_vector(0 downto 0);
    writeModule1_call_data : out  std_logic_vector(103 downto 0);
    writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
    writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_return_acks : in   std_logic_vector(0 downto 0);
    writeModule1_return_data : in   std_logic_vector(0 downto 0);
    writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ct_core;
architecture ct_core_arch of ct_core is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 176)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal inp_d0_buffer :  std_logic_vector(15 downto 0);
  signal inp_d0_update_enable: Boolean;
  signal inp_d1_buffer :  std_logic_vector(15 downto 0);
  signal inp_d1_update_enable: Boolean;
  signal inp_d2_buffer :  std_logic_vector(15 downto 0);
  signal inp_d2_update_enable: Boolean;
  signal ker_d1_buffer :  std_logic_vector(15 downto 0);
  signal ker_d1_update_enable: Boolean;
  signal ker_d2_buffer :  std_logic_vector(15 downto 0);
  signal ker_d2_update_enable: Boolean;
  signal out_d0_buffer :  std_logic_vector(15 downto 0);
  signal out_d0_update_enable: Boolean;
  signal out_d1_buffer :  std_logic_vector(15 downto 0);
  signal out_d1_update_enable: Boolean;
  signal out_d2_buffer :  std_logic_vector(15 downto 0);
  signal out_d2_update_enable: Boolean;
  signal stride_buffer :  std_logic_vector(15 downto 0);
  signal stride_update_enable: Boolean;
  signal padding_buffer :  std_logic_vector(15 downto 0);
  signal padding_update_enable: Boolean;
  signal index1_buffer :  std_logic_vector(7 downto 0);
  signal index1_update_enable: Boolean;
  signal index3_buffer :  std_logic_vector(7 downto 0);
  signal index3_update_enable: Boolean;
  -- output port buffer signals
  signal ct_core_CP_345_start: Boolean;
  signal ct_core_CP_345_symbol: Boolean;
  -- volatile/operator module components. 
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal phi_stmt_132_ack_0 : boolean;
  signal W_dim2_limit_180_delayed_1_0_181_inst_ack_1 : boolean;
  signal phi_stmt_132_req_1 : boolean;
  signal next_add_dest_dim1_262_131_buf_req_1 : boolean;
  signal SUB_u16_u16_294_inst_req_1 : boolean;
  signal W_dim2_limit_180_delayed_1_0_181_inst_req_1 : boolean;
  signal call_stmt_166_call_ack_0 : boolean;
  signal call_stmt_166_call_req_0 : boolean;
  signal next_add_dest_dim0_268_127_buf_ack_1 : boolean;
  signal next_add_dest_dim0_268_127_buf_req_1 : boolean;
  signal add_dest_dim1_init_105_130_buf_ack_0 : boolean;
  signal W_nid1_true3_233_delayed_1_0_240_inst_ack_1 : boolean;
  signal next_add_dest_dim0_268_127_buf_ack_0 : boolean;
  signal next_add_dest_dim1_262_131_buf_ack_0 : boolean;
  signal next_add_dest_dim0_268_127_buf_req_0 : boolean;
  signal next_add_dest_dim1_262_131_buf_req_0 : boolean;
  signal type_cast_169_inst_ack_1 : boolean;
  signal add_dest_dim1_init_105_130_buf_req_0 : boolean;
  signal next_add_src_252_135_buf_ack_0 : boolean;
  signal type_cast_169_inst_req_1 : boolean;
  signal do_while_stmt_110_branch_ack_0 : boolean;
  signal call_stmt_175_call_ack_1 : boolean;
  signal phi_stmt_112_ack_0 : boolean;
  signal add_dest_dim0_init_100_126_buf_ack_0 : boolean;
  signal SUB_u16_u16_192_inst_ack_1 : boolean;
  signal SUB_u16_u16_192_inst_req_1 : boolean;
  signal W_dim2_limit_180_delayed_1_0_181_inst_ack_0 : boolean;
  signal call_stmt_175_call_req_1 : boolean;
  signal add_dest_dim1_init_105_130_buf_ack_1 : boolean;
  signal phi_stmt_132_req_0 : boolean;
  signal W_dim2_limit_180_delayed_1_0_181_inst_req_0 : boolean;
  signal W_nid1_true3_233_delayed_1_0_240_inst_req_1 : boolean;
  signal SUB_u16_u16_192_inst_ack_0 : boolean;
  signal SUB_u16_u16_192_inst_req_0 : boolean;
  signal next_add_src_252_135_buf_req_0 : boolean;
  signal add_dest_dim1_init_105_130_buf_req_1 : boolean;
  signal type_cast_169_inst_ack_0 : boolean;
  signal phi_stmt_128_req_1 : boolean;
  signal SUB_u16_u16_294_inst_req_0 : boolean;
  signal SUB_u16_u16_294_inst_ack_1 : boolean;
  signal do_while_stmt_110_branch_ack_1 : boolean;
  signal call_stmt_166_call_ack_1 : boolean;
  signal add_dest_dim0_init_100_126_buf_ack_1 : boolean;
  signal W_nid1_true3_233_delayed_1_0_240_inst_ack_0 : boolean;
  signal call_stmt_175_call_ack_0 : boolean;
  signal type_cast_169_inst_req_0 : boolean;
  signal add_dest_dim0_init_100_126_buf_req_1 : boolean;
  signal do_while_stmt_110_branch_req_0 : boolean;
  signal call_stmt_166_call_req_1 : boolean;
  signal call_stmt_175_call_req_0 : boolean;
  signal phi_stmt_112_req_1 : boolean;
  signal phi_stmt_112_req_0 : boolean;
  signal next_input_dim0_290_115_buf_req_0 : boolean;
  signal next_input_dim0_290_115_buf_ack_0 : boolean;
  signal next_input_dim0_290_115_buf_req_1 : boolean;
  signal next_input_dim0_290_115_buf_ack_1 : boolean;
  signal W_nid1_true3_233_delayed_1_0_240_inst_req_0 : boolean;
  signal SUB_u16_u16_294_inst_ack_0 : boolean;
  signal phi_stmt_116_req_1 : boolean;
  signal phi_stmt_116_req_0 : boolean;
  signal phi_stmt_116_ack_0 : boolean;
  signal next_add_dest_dim1_262_131_buf_ack_1 : boolean;
  signal next_input_dim1_284_119_buf_req_0 : boolean;
  signal next_input_dim1_284_119_buf_ack_0 : boolean;
  signal next_input_dim1_284_119_buf_req_1 : boolean;
  signal next_input_dim1_284_119_buf_ack_1 : boolean;
  signal add_dest_dim0_init_100_126_buf_req_0 : boolean;
  signal phi_stmt_128_ack_0 : boolean;
  signal phi_stmt_120_req_1 : boolean;
  signal phi_stmt_120_req_0 : boolean;
  signal next_add_src_252_135_buf_ack_1 : boolean;
  signal phi_stmt_120_ack_0 : boolean;
  signal next_add_src_252_135_buf_req_1 : boolean;
  signal phi_stmt_128_req_0 : boolean;
  signal next_input_dim2_274_123_buf_req_0 : boolean;
  signal next_input_dim2_274_123_buf_ack_0 : boolean;
  signal next_input_dim2_274_123_buf_req_1 : boolean;
  signal next_input_dim2_274_123_buf_ack_1 : boolean;
  signal phi_stmt_124_req_1 : boolean;
  signal phi_stmt_124_req_0 : boolean;
  signal phi_stmt_124_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ct_core_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 176) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= inp_d0;
  inp_d0_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= inp_d1;
  inp_d1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= inp_d2;
  inp_d2_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= ker_d1;
  ker_d1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= ker_d2;
  ker_d2_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= out_d0;
  out_d0_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(111 downto 96) <= out_d1;
  out_d1_buffer <= in_buffer_data_out(111 downto 96);
  in_buffer_data_in(127 downto 112) <= out_d2;
  out_d2_buffer <= in_buffer_data_out(127 downto 112);
  in_buffer_data_in(143 downto 128) <= stride;
  stride_buffer <= in_buffer_data_out(143 downto 128);
  in_buffer_data_in(159 downto 144) <= padding;
  padding_buffer <= in_buffer_data_out(159 downto 144);
  in_buffer_data_in(167 downto 160) <= index1;
  index1_buffer <= in_buffer_data_out(167 downto 160);
  in_buffer_data_in(175 downto 168) <= index3;
  index3_buffer <= in_buffer_data_out(175 downto 168);
  in_buffer_data_in(tag_length + 175 downto 176) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 175 downto 176);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ct_core_CP_345_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ct_core_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ct_core_CP_345_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ct_core_CP_345_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ct_core_CP_345_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ct_core_CP_345: Block -- control-path 
    signal ct_core_CP_345_elements: BooleanArray(159 downto 0);
    -- 
  begin -- 
    ct_core_CP_345_elements(0) <= ct_core_CP_345_start;
    ct_core_CP_345_symbol <= ct_core_CP_345_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_78/$entry
      -- CP-element group 0: 	 branch_block_stmt_78/branch_block_stmt_78__entry__
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_82_to_assign_stmt_109__entry__
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_82_to_assign_stmt_109__exit__
      -- CP-element group 0: 	 branch_block_stmt_78/do_while_stmt_110__entry__
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_82_to_assign_stmt_109/$entry
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_82_to_assign_stmt_109/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	159 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_78/$exit
      -- CP-element group 1: 	 branch_block_stmt_78/branch_block_stmt_78__exit__
      -- CP-element group 1: 	 branch_block_stmt_78/do_while_stmt_110__exit__
      -- 
    ct_core_CP_345_elements(1) <= ct_core_CP_345_elements(159);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_78/do_while_stmt_110/$entry
      -- CP-element group 2: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110__entry__
      -- 
    ct_core_CP_345_elements(2) <= ct_core_CP_345_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	159 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110__exit__
      -- 
    -- Element group ct_core_CP_345_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_78/do_while_stmt_110/loop_back
      -- 
    -- Element group ct_core_CP_345_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	157 
    -- CP-element group 5: 	158 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_78/do_while_stmt_110/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_78/do_while_stmt_110/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_78/do_while_stmt_110/condition_done
      -- 
    ct_core_CP_345_elements(5) <= ct_core_CP_345_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	156 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_78/do_while_stmt_110/loop_body_done
      -- 
    ct_core_CP_345_elements(6) <= ct_core_CP_345_elements(156);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	114 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	95 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/back_edge_to_loop_body
      -- 
    ct_core_CP_345_elements(7) <= ct_core_CP_345_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	116 
    -- CP-element group 8: 	97 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	78 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/first_time_through_loop_body
      -- 
    ct_core_CP_345_elements(8) <= ct_core_CP_345_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	109 
    -- CP-element group 9: 	143 
    -- CP-element group 9: 	147 
    -- CP-element group 9: 	139 
    -- CP-element group 9: 	151 
    -- CP-element group 9: 	155 
    -- CP-element group 9: 	108 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	90 
    -- CP-element group 9: 	89 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	70 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/loop_body_start
      -- 
    -- Element group ct_core_CP_345_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	142 
    -- CP-element group 10: 	146 
    -- CP-element group 10: 	154 
    -- CP-element group 10: 	155 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/condition_evaluated
      -- 
    condition_evaluated_374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(10), ack => do_while_stmt_110_branch_req_0); -- 
    ct_core_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(142) & ct_core_CP_345_elements(146) & ct_core_CP_345_elements(154) & ct_core_CP_345_elements(155) & ct_core_CP_345_elements(14);
      gj_ct_core_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	108 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	89 
    -- CP-element group 11: 	70 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	110 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	72 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_sample_start__ps
      -- 
    ct_core_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(34) & ct_core_CP_345_elements(51) & ct_core_CP_345_elements(108) & ct_core_CP_345_elements(15) & ct_core_CP_345_elements(89) & ct_core_CP_345_elements(70) & ct_core_CP_345_elements(14);
      gj_ct_core_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	111 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	92 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	144 
    -- CP-element group 12: 	148 
    -- CP-element group 12: 	140 
    -- CP-element group 12: 	156 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	108 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	89 
    -- CP-element group 12: 	70 
    -- CP-element group 12:  members (7) 
      -- CP-element group 12: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_sample_completed_
      -- 
    ct_core_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(36) & ct_core_CP_345_elements(54) & ct_core_CP_345_elements(111) & ct_core_CP_345_elements(18) & ct_core_CP_345_elements(73) & ct_core_CP_345_elements(92);
      gj_ct_core_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	109 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	90 
    -- CP-element group 13: 	71 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	112 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	93 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_update_start__ps
      -- 
    ct_core_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(35) & ct_core_CP_345_elements(52) & ct_core_CP_345_elements(109) & ct_core_CP_345_elements(16) & ct_core_CP_345_elements(90) & ct_core_CP_345_elements(71);
      gj_ct_core_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	113 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	94 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/aggregated_phi_update_ack
      -- 
    ct_core_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(37) & ct_core_CP_345_elements(56) & ct_core_CP_345_elements(113) & ct_core_CP_345_elements(20) & ct_core_CP_345_elements(75) & ct_core_CP_345_elements(94);
      gj_ct_core_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	142 
    -- CP-element group 15: 	146 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_sample_start_
      -- 
    ct_core_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(142) & ct_core_CP_345_elements(146) & ct_core_CP_345_elements(12);
      gj_ct_core_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_update_start_
      -- 
    ct_core_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(20);
      gj_ct_core_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_sample_start__ps
      -- 
    ct_core_CP_345_elements(17) <= ct_core_CP_345_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_sample_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_update_start__ps
      -- 
    ct_core_CP_345_elements(19) <= ct_core_CP_345_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_update_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_loopback_trigger
      -- 
    ct_core_CP_345_elements(21) <= ct_core_CP_345_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_loopback_sample_req_ps
      -- 
    phi_stmt_112_loopback_sample_req_389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_loopback_sample_req_389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(22), ack => phi_stmt_112_req_1); -- 
    -- Element group ct_core_CP_345_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_entry_trigger
      -- 
    ct_core_CP_345_elements(23) <= ct_core_CP_345_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_entry_sample_req_ps
      -- 
    phi_stmt_112_entry_sample_req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_entry_sample_req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(24), ack => phi_stmt_112_req_0); -- 
    -- Element group ct_core_CP_345_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_112_phi_mux_ack_ps
      -- 
    phi_stmt_112_phi_mux_ack_395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_112_ack_0, ack => ct_core_CP_345_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_sample_completed_
      -- 
    -- Element group ct_core_CP_345_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_update_start_
      -- 
    -- Element group ct_core_CP_345_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_update_completed__ps
      -- 
    ct_core_CP_345_elements(28) <= ct_core_CP_345_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim0_init_114_update_completed_
      -- 
    -- Element group ct_core_CP_345_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => ct_core_CP_345_elements(27), ack => ct_core_CP_345_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Sample/req
      -- 
    req_416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(30), ack => next_input_dim0_290_115_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_update_start_
      -- CP-element group 31: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Update/req
      -- 
    req_421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(31), ack => next_input_dim0_290_115_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Sample/ack
      -- 
    ack_417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_290_115_buf_ack_0, ack => ct_core_CP_345_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim0_115_Update/ack
      -- 
    ack_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_290_115_buf_ack_1, ack => ct_core_CP_345_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	142 
    -- CP-element group 34: 	146 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_sample_start_
      -- 
    ct_core_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(142) & ct_core_CP_345_elements(146) & ct_core_CP_345_elements(12);
      gj_ct_core_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_update_start_
      -- 
    ct_core_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(37);
      gj_ct_core_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	12 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_sample_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(36) is bound as output of CP function.
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_update_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_loopback_trigger
      -- 
    ct_core_CP_345_elements(38) <= ct_core_CP_345_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_loopback_sample_req_ps
      -- 
    phi_stmt_116_loopback_sample_req_433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_loopback_sample_req_433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(39), ack => phi_stmt_116_req_1); -- 
    -- Element group ct_core_CP_345_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_entry_trigger
      -- 
    ct_core_CP_345_elements(40) <= ct_core_CP_345_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_entry_sample_req_ps
      -- 
    phi_stmt_116_entry_sample_req_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_entry_sample_req_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(41), ack => phi_stmt_116_req_0); -- 
    -- Element group ct_core_CP_345_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_116_phi_mux_ack_ps
      -- 
    phi_stmt_116_phi_mux_ack_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_116_ack_0, ack => ct_core_CP_345_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_sample_completed_
      -- 
    -- Element group ct_core_CP_345_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_update_start_
      -- 
    -- Element group ct_core_CP_345_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_update_completed__ps
      -- 
    ct_core_CP_345_elements(45) <= ct_core_CP_345_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim1_init_118_update_completed_
      -- 
    -- Element group ct_core_CP_345_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => ct_core_CP_345_elements(44), ack => ct_core_CP_345_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Sample/req
      -- 
    req_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(47), ack => next_input_dim1_284_119_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_update_start_
      -- CP-element group 48: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Update/req
      -- 
    req_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(48), ack => next_input_dim1_284_119_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Sample/ack
      -- 
    ack_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_284_119_buf_ack_0, ack => ct_core_CP_345_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim1_119_Update/ack
      -- 
    ack_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_284_119_buf_ack_1, ack => ct_core_CP_345_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	142 
    -- CP-element group 51: 	12 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_sample_start_
      -- 
    ct_core_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(142) & ct_core_CP_345_elements(12);
      gj_ct_core_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	133 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_update_start_
      -- 
    ct_core_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(133);
      gj_ct_core_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_sample_start__ps
      -- 
    ct_core_CP_345_elements(53) <= ct_core_CP_345_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_sample_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_update_start__ps
      -- 
    ct_core_CP_345_elements(55) <= ct_core_CP_345_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	131 
    -- CP-element group 56: 	14 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_update_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_loopback_trigger
      -- 
    ct_core_CP_345_elements(57) <= ct_core_CP_345_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_loopback_sample_req_ps
      -- 
    phi_stmt_120_loopback_sample_req_477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_120_loopback_sample_req_477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(58), ack => phi_stmt_120_req_1); -- 
    -- Element group ct_core_CP_345_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_entry_trigger
      -- 
    ct_core_CP_345_elements(59) <= ct_core_CP_345_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_entry_sample_req_ps
      -- 
    phi_stmt_120_entry_sample_req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_120_entry_sample_req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(60), ack => phi_stmt_120_req_0); -- 
    -- Element group ct_core_CP_345_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_120_phi_mux_ack_ps
      -- 
    phi_stmt_120_phi_mux_ack_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_120_ack_0, ack => ct_core_CP_345_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_sample_completed_
      -- 
    -- Element group ct_core_CP_345_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_update_start_
      -- 
    -- Element group ct_core_CP_345_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_update_completed__ps
      -- 
    ct_core_CP_345_elements(64) <= ct_core_CP_345_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_input_dim2_init_122_update_completed_
      -- 
    -- Element group ct_core_CP_345_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => ct_core_CP_345_elements(63), ack => ct_core_CP_345_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Sample/req
      -- 
    req_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(66), ack => next_input_dim2_274_123_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_update_start_
      -- CP-element group 67: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Update/req
      -- 
    req_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(67), ack => next_input_dim2_274_123_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Sample/ack
      -- 
    ack_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_274_123_buf_ack_0, ack => ct_core_CP_345_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_input_dim2_123_Update/ack
      -- 
    ack_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_274_123_buf_ack_1, ack => ct_core_CP_345_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	142 
    -- CP-element group 70: 	146 
    -- CP-element group 70: 	12 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_sample_start_
      -- 
    ct_core_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(142) & ct_core_CP_345_elements(146) & ct_core_CP_345_elements(12);
      gj_ct_core_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	133 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_update_start_
      -- 
    ct_core_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(133);
      gj_ct_core_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_sample_start__ps
      -- 
    ct_core_CP_345_elements(72) <= ct_core_CP_345_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_sample_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_update_start__ps
      -- 
    ct_core_CP_345_elements(74) <= ct_core_CP_345_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	131 
    -- CP-element group 75: 	14 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_update_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_loopback_trigger
      -- 
    ct_core_CP_345_elements(76) <= ct_core_CP_345_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_loopback_sample_req_ps
      -- 
    phi_stmt_124_loopback_sample_req_521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_loopback_sample_req_521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(77), ack => phi_stmt_124_req_1); -- 
    -- Element group ct_core_CP_345_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_entry_trigger
      -- 
    ct_core_CP_345_elements(78) <= ct_core_CP_345_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_entry_sample_req_ps
      -- 
    phi_stmt_124_entry_sample_req_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_entry_sample_req_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(79), ack => phi_stmt_124_req_0); -- 
    -- Element group ct_core_CP_345_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_phi_mux_ack_ps
      -- CP-element group 80: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_124_phi_mux_ack
      -- 
    phi_stmt_124_phi_mux_ack_527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_124_ack_0, ack => ct_core_CP_345_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Sample/req
      -- 
    req_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(81), ack => add_dest_dim0_init_100_126_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_update_start_
      -- CP-element group 82: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Update/req
      -- CP-element group 82: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Update/$entry
      -- 
    req_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(82), ack => add_dest_dim0_init_100_126_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_sample_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Sample/ack
      -- CP-element group 83: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_sample_completed_
      -- 
    ack_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_100_126_buf_ack_0, ack => ct_core_CP_345_elements(83)); -- 
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_update_completed__ps
      -- CP-element group 84: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Update/ack
      -- CP-element group 84: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim0_init_126_Update/$exit
      -- 
    ack_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_100_126_buf_ack_1, ack => ct_core_CP_345_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_sample_start__ps
      -- 
    req_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(85), ack => next_add_dest_dim0_268_127_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Update/req
      -- CP-element group 86: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_update_start_
      -- CP-element group 86: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_update_start__ps
      -- 
    req_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(86), ack => next_add_dest_dim0_268_127_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_sample_completed__ps
      -- 
    ack_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_268_127_buf_ack_0, ack => ct_core_CP_345_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim0_127_update_completed__ps
      -- 
    ack_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_268_127_buf_ack_1, ack => ct_core_CP_345_elements(88)); -- 
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	9 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	142 
    -- CP-element group 89: 	146 
    -- CP-element group 89: 	150 
    -- CP-element group 89: 	12 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	11 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_sample_start_
      -- 
    ct_core_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(142) & ct_core_CP_345_elements(146) & ct_core_CP_345_elements(150) & ct_core_CP_345_elements(12);
      gj_ct_core_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	9 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	133 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	13 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_update_start_
      -- 
    ct_core_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(133);
      gj_ct_core_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	11 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_sample_start__ps
      -- 
    ct_core_CP_345_elements(91) <= ct_core_CP_345_elements(11);
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	12 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_sample_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(92) is bound as output of CP function.
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	13 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_update_start__ps
      -- 
    ct_core_CP_345_elements(93) <= ct_core_CP_345_elements(13);
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	131 
    -- CP-element group 94: 	14 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_update_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	7 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_loopback_trigger
      -- 
    ct_core_CP_345_elements(95) <= ct_core_CP_345_elements(7);
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_loopback_sample_req_ps
      -- CP-element group 96: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_loopback_sample_req
      -- 
    phi_stmt_128_loopback_sample_req_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_128_loopback_sample_req_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(96), ack => phi_stmt_128_req_1); -- 
    -- Element group ct_core_CP_345_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	8 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_entry_trigger
      -- 
    ct_core_CP_345_elements(97) <= ct_core_CP_345_elements(8);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_entry_sample_req_ps
      -- CP-element group 98: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_entry_sample_req
      -- 
    phi_stmt_128_entry_sample_req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_128_entry_sample_req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(98), ack => phi_stmt_128_req_0); -- 
    -- Element group ct_core_CP_345_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_phi_mux_ack_ps
      -- CP-element group 99: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_128_phi_mux_ack
      -- 
    phi_stmt_128_phi_mux_ack_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_128_ack_0, ack => ct_core_CP_345_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Sample/req
      -- CP-element group 100: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_sample_start__ps
      -- 
    req_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(100), ack => add_dest_dim1_init_105_130_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_update_start_
      -- CP-element group 101: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Update/req
      -- CP-element group 101: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_update_start__ps
      -- 
    req_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(101), ack => add_dest_dim1_init_105_130_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Sample/ack
      -- CP-element group 102: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_sample_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_sample_completed_
      -- 
    ack_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_105_130_buf_ack_0, ack => ct_core_CP_345_elements(102)); -- 
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Update/ack
      -- CP-element group 103: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_update_completed__ps
      -- CP-element group 103: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_dest_dim1_init_130_Update/$exit
      -- 
    ack_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_105_130_buf_ack_1, ack => ct_core_CP_345_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Sample/req
      -- CP-element group 104: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_sample_start__ps
      -- 
    req_612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(104), ack => next_add_dest_dim1_262_131_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Update/req
      -- CP-element group 105: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_update_start_
      -- CP-element group 105: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_update_start__ps
      -- 
    req_617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(105), ack => next_add_dest_dim1_262_131_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Sample/ack
      -- CP-element group 106: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_sample_completed__ps
      -- 
    ack_613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_262_131_buf_ack_0, ack => ct_core_CP_345_elements(106)); -- 
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_dest_dim1_131_Update/ack
      -- 
    ack_618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_262_131_buf_ack_1, ack => ct_core_CP_345_elements(107)); -- 
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	9 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	12 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	11 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_sample_start_
      -- 
    ct_core_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(12);
      gj_ct_core_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	9 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	129 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	13 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_update_start_
      -- 
    ct_core_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(129);
      gj_ct_core_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	11 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_sample_start__ps
      -- 
    ct_core_CP_345_elements(110) <= ct_core_CP_345_elements(11);
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	12 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_sample_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(111) is bound as output of CP function.
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	13 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_update_start__ps
      -- 
    ct_core_CP_345_elements(112) <= ct_core_CP_345_elements(13);
    -- CP-element group 113:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	127 
    -- CP-element group 113: 	14 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_update_completed_
      -- 
    -- Element group ct_core_CP_345_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	7 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_loopback_trigger
      -- 
    ct_core_CP_345_elements(114) <= ct_core_CP_345_elements(7);
    -- CP-element group 115:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_loopback_sample_req
      -- CP-element group 115: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_loopback_sample_req_ps
      -- 
    phi_stmt_132_loopback_sample_req_629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_132_loopback_sample_req_629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(115), ack => phi_stmt_132_req_1); -- 
    -- Element group ct_core_CP_345_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	8 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_entry_trigger
      -- 
    ct_core_CP_345_elements(116) <= ct_core_CP_345_elements(8);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_entry_sample_req_ps
      -- CP-element group 117: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_entry_sample_req
      -- 
    phi_stmt_132_entry_sample_req_632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_132_entry_sample_req_632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(117), ack => phi_stmt_132_req_0); -- 
    -- Element group ct_core_CP_345_elements(117) is bound as output of CP function.
    -- CP-element group 118:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_phi_mux_ack
      -- CP-element group 118: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/phi_stmt_132_phi_mux_ack_ps
      -- 
    phi_stmt_132_phi_mux_ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_132_ack_0, ack => ct_core_CP_345_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_sample_start__ps
      -- CP-element group 119: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_sample_completed__ps
      -- 
    -- Element group ct_core_CP_345_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_update_start_
      -- CP-element group 120: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_update_start__ps
      -- 
    -- Element group ct_core_CP_345_elements(120) is bound as output of CP function.
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_update_completed__ps
      -- 
    ct_core_CP_345_elements(121) <= ct_core_CP_345_elements(122);
    -- CP-element group 122:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	121 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_add_src_init_134_update_completed_
      -- 
    -- Element group ct_core_CP_345_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => ct_core_CP_345_elements(120), ack => ct_core_CP_345_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_sample_start__ps
      -- CP-element group 123: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Sample/req
      -- CP-element group 123: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_sample_start_
      -- 
    req_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(123), ack => next_add_src_252_135_buf_req_0); -- 
    -- Element group ct_core_CP_345_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_update_start_
      -- CP-element group 124: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_update_start__ps
      -- CP-element group 124: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Update/req
      -- 
    req_661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(124), ack => next_add_src_252_135_buf_req_1); -- 
    -- Element group ct_core_CP_345_elements(124) is bound as output of CP function.
    -- CP-element group 125:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Sample/ack
      -- CP-element group 125: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_sample_completed__ps
      -- 
    ack_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_252_135_buf_ack_0, ack => ct_core_CP_345_elements(125)); -- 
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_update_completed__ps
      -- CP-element group 126: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/R_next_add_src_135_Update/ack
      -- 
    ack_662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_252_135_buf_ack_1, ack => ct_core_CP_345_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	113 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Sample/crr
      -- CP-element group 127: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_sample_start_
      -- 
    crr_671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(127), ack => call_stmt_166_call_req_0); -- 
    ct_core_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(113) & ct_core_CP_345_elements(129);
      gj_ct_core_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	137 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_update_start_
      -- CP-element group 128: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Update/ccr
      -- 
    ccr_676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(128), ack => call_stmt_166_call_req_1); -- 
    ct_core_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ct_core_CP_345_elements(137);
      gj_ct_core_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	109 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Sample/cra
      -- CP-element group 129: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_sample_completed_
      -- 
    cra_672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_166_call_ack_0, ack => ct_core_CP_345_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	135 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Update/cca
      -- CP-element group 130: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_166_Update/$exit
      -- 
    cca_677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_166_call_ack_1, ack => ct_core_CP_345_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	56 
    -- CP-element group 131: 	75 
    -- CP-element group 131: 	94 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Sample/rr
      -- 
    rr_685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(131), ack => type_cast_169_inst_req_0); -- 
    ct_core_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(56) & ct_core_CP_345_elements(75) & ct_core_CP_345_elements(94) & ct_core_CP_345_elements(133);
      gj_ct_core_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	137 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_update_start_
      -- 
    cr_690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(132), ack => type_cast_169_inst_req_1); -- 
    ct_core_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ct_core_CP_345_elements(137);
      gj_ct_core_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	52 
    -- CP-element group 133: 	131 
    -- CP-element group 133: 	90 
    -- CP-element group 133: 	71 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_sample_completed_
      -- 
    ra_686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_0, ack => ct_core_CP_345_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/type_cast_169_update_completed_
      -- 
    ca_691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_1, ack => ct_core_CP_345_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: 	130 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Sample/crr
      -- 
    crr_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(135), ack => call_stmt_175_call_req_0); -- 
    ct_core_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(134) & ct_core_CP_345_elements(130) & ct_core_CP_345_elements(137);
      gj_ct_core_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_update_start_
      -- CP-element group 136: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Update/ccr
      -- CP-element group 136: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Update/$entry
      -- 
    ccr_704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(136), ack => call_stmt_175_call_req_1); -- 
    ct_core_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ct_core_CP_345_elements(138);
      gj_ct_core_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: 	128 
    -- CP-element group 137: 	132 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Sample/cra
      -- CP-element group 137: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Sample/$exit
      -- 
    cra_700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_175_call_ack_0, ack => ct_core_CP_345_elements(137)); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	156 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Update/cca
      -- CP-element group 138: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/call_stmt_175_Update/$exit
      -- 
    cca_705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_175_call_ack_1, ack => ct_core_CP_345_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	9 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Sample/req
      -- CP-element group 139: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Sample/$entry
      -- 
    req_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(139), ack => W_dim2_limit_180_delayed_1_0_181_inst_req_0); -- 
    ct_core_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(141);
      gj_ct_core_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	12 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Update/req
      -- CP-element group 140: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_update_start_
      -- 
    req_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(140), ack => W_dim2_limit_180_delayed_1_0_181_inst_req_1); -- 
    ct_core_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(12) & ct_core_CP_345_elements(142);
      gj_ct_core_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Sample/ack
      -- CP-element group 141: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Sample/$exit
      -- 
    ack_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_180_delayed_1_0_181_inst_ack_0, ack => ct_core_CP_345_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	10 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	34 
    -- CP-element group 142: 	51 
    -- CP-element group 142: 	140 
    -- CP-element group 142: 	15 
    -- CP-element group 142: 	89 
    -- CP-element group 142: 	70 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Update/ack
      -- CP-element group 142: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_183_update_completed_
      -- 
    ack_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_180_delayed_1_0_181_inst_ack_1, ack => ct_core_CP_345_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	9 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_sample_start_
      -- 
    rr_727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(143), ack => SUB_u16_u16_192_inst_req_0); -- 
    ct_core_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(145);
      gj_ct_core_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	12 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_update_start_
      -- 
    cr_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(144), ack => SUB_u16_u16_192_inst_req_1); -- 
    ct_core_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(12) & ct_core_CP_345_elements(146);
      gj_ct_core_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_sample_completed_
      -- 
    ra_728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_192_inst_ack_0, ack => ct_core_CP_345_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	10 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	34 
    -- CP-element group 146: 	144 
    -- CP-element group 146: 	15 
    -- CP-element group 146: 	89 
    -- CP-element group 146: 	70 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_192_update_completed_
      -- 
    ca_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_192_inst_ack_1, ack => ct_core_CP_345_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	9 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Sample/req
      -- 
    req_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(147), ack => W_nid1_true3_233_delayed_1_0_240_inst_req_0); -- 
    ct_core_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(149);
      gj_ct_core_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	12 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_update_start_
      -- CP-element group 148: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Update/req
      -- CP-element group 148: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Update/$entry
      -- 
    req_746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(148), ack => W_nid1_true3_233_delayed_1_0_240_inst_req_1); -- 
    ct_core_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(12) & ct_core_CP_345_elements(150);
      gj_ct_core_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Sample/ack
      -- CP-element group 149: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Sample/$exit
      -- 
    ack_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true3_233_delayed_1_0_240_inst_ack_0, ack => ct_core_CP_345_elements(149)); -- 
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	156 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: 	89 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Update/ack
      -- CP-element group 150: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/assign_stmt_242_Update/$exit
      -- 
    ack_747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true3_233_delayed_1_0_240_inst_ack_1, ack => ct_core_CP_345_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	9 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_sample_start_
      -- 
    rr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(151), ack => SUB_u16_u16_294_inst_req_0); -- 
    ct_core_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(9) & ct_core_CP_345_elements(153);
      gj_ct_core_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Update/cr
      -- CP-element group 152: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_update_start_
      -- 
    cr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_345_elements(152), ack => SUB_u16_u16_294_inst_req_1); -- 
    ct_core_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ct_core_CP_345_elements(154);
      gj_ct_core_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Sample/ra
      -- 
    ra_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_294_inst_ack_0, ack => ct_core_CP_345_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	10 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/SUB_u16_u16_294_Update/ca
      -- 
    ca_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_294_inst_ack_1, ack => ct_core_CP_345_elements(154)); -- 
    -- CP-element group 155:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	9 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	10 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group ct_core_CP_345_elements(155) is a control-delay.
    cp_element_155_delay: control_delay_element  generic map(name => " 155_delay", delay_value => 1)  port map(req => ct_core_CP_345_elements(9), ack => ct_core_CP_345_elements(155), clk => clk, reset =>reset);
    -- CP-element group 156:  join  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	138 
    -- CP-element group 156: 	150 
    -- CP-element group 156: 	12 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	6 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_78/do_while_stmt_110/do_while_stmt_110_loop_body/$exit
      -- 
    ct_core_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_345_elements(138) & ct_core_CP_345_elements(150) & ct_core_CP_345_elements(12);
      gj_ct_core_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_345_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	5 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (2) 
      -- CP-element group 157: 	 branch_block_stmt_78/do_while_stmt_110/loop_exit/$exit
      -- CP-element group 157: 	 branch_block_stmt_78/do_while_stmt_110/loop_exit/ack
      -- 
    ack_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_110_branch_ack_0, ack => ct_core_CP_345_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	5 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_78/do_while_stmt_110/loop_taken/$exit
      -- CP-element group 158: 	 branch_block_stmt_78/do_while_stmt_110/loop_taken/ack
      -- 
    ack_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_110_branch_ack_1, ack => ct_core_CP_345_elements(158)); -- 
    -- CP-element group 159:  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	3 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	1 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_78/do_while_stmt_110/$exit
      -- 
    ct_core_CP_345_elements(159) <= ct_core_CP_345_elements(3);
    ct_core_do_while_stmt_110_terminator_771: loop_terminator -- 
      generic map (name => " ct_core_do_while_stmt_110_terminator_771", max_iterations_in_flight =>15) 
      port map(loop_body_exit => ct_core_CP_345_elements(6),loop_continue => ct_core_CP_345_elements(158),loop_terminate => ct_core_CP_345_elements(157),loop_back => ct_core_CP_345_elements(4),loop_exit => ct_core_CP_345_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_112_phi_seq_423_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_345_elements(23);
      ct_core_CP_345_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_345_elements(26);
      ct_core_CP_345_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_345_elements(28);
      ct_core_CP_345_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_345_elements(21);
      ct_core_CP_345_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_345_elements(32);
      ct_core_CP_345_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_345_elements(33);
      ct_core_CP_345_elements(22) <= phi_mux_reqs(1);
      phi_stmt_112_phi_seq_423 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_112_phi_seq_423") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_345_elements(17), 
          phi_sample_ack => ct_core_CP_345_elements(18), 
          phi_update_req => ct_core_CP_345_elements(19), 
          phi_update_ack => ct_core_CP_345_elements(20), 
          phi_mux_ack => ct_core_CP_345_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_116_phi_seq_467_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_345_elements(40);
      ct_core_CP_345_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_345_elements(43);
      ct_core_CP_345_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_345_elements(45);
      ct_core_CP_345_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_345_elements(38);
      ct_core_CP_345_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_345_elements(49);
      ct_core_CP_345_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_345_elements(50);
      ct_core_CP_345_elements(39) <= phi_mux_reqs(1);
      phi_stmt_116_phi_seq_467 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_116_phi_seq_467") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_345_elements(11), 
          phi_sample_ack => ct_core_CP_345_elements(36), 
          phi_update_req => ct_core_CP_345_elements(13), 
          phi_update_ack => ct_core_CP_345_elements(37), 
          phi_mux_ack => ct_core_CP_345_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_120_phi_seq_511_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_345_elements(59);
      ct_core_CP_345_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_345_elements(62);
      ct_core_CP_345_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_345_elements(64);
      ct_core_CP_345_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_345_elements(57);
      ct_core_CP_345_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_345_elements(68);
      ct_core_CP_345_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_345_elements(69);
      ct_core_CP_345_elements(58) <= phi_mux_reqs(1);
      phi_stmt_120_phi_seq_511 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_120_phi_seq_511") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_345_elements(53), 
          phi_sample_ack => ct_core_CP_345_elements(54), 
          phi_update_req => ct_core_CP_345_elements(55), 
          phi_update_ack => ct_core_CP_345_elements(56), 
          phi_mux_ack => ct_core_CP_345_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_124_phi_seq_565_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_345_elements(78);
      ct_core_CP_345_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_345_elements(83);
      ct_core_CP_345_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_345_elements(84);
      ct_core_CP_345_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_345_elements(76);
      ct_core_CP_345_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_345_elements(87);
      ct_core_CP_345_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_345_elements(88);
      ct_core_CP_345_elements(77) <= phi_mux_reqs(1);
      phi_stmt_124_phi_seq_565 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_124_phi_seq_565") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_345_elements(72), 
          phi_sample_ack => ct_core_CP_345_elements(73), 
          phi_update_req => ct_core_CP_345_elements(74), 
          phi_update_ack => ct_core_CP_345_elements(75), 
          phi_mux_ack => ct_core_CP_345_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_128_phi_seq_619_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_345_elements(97);
      ct_core_CP_345_elements(100)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_345_elements(102);
      ct_core_CP_345_elements(101)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_345_elements(103);
      ct_core_CP_345_elements(98) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_345_elements(95);
      ct_core_CP_345_elements(104)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_345_elements(106);
      ct_core_CP_345_elements(105)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_345_elements(107);
      ct_core_CP_345_elements(96) <= phi_mux_reqs(1);
      phi_stmt_128_phi_seq_619 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_128_phi_seq_619") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_345_elements(91), 
          phi_sample_ack => ct_core_CP_345_elements(92), 
          phi_update_req => ct_core_CP_345_elements(93), 
          phi_update_ack => ct_core_CP_345_elements(94), 
          phi_mux_ack => ct_core_CP_345_elements(99), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_132_phi_seq_663_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_345_elements(116);
      ct_core_CP_345_elements(119)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_345_elements(119);
      ct_core_CP_345_elements(120)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_345_elements(121);
      ct_core_CP_345_elements(117) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_345_elements(114);
      ct_core_CP_345_elements(123)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_345_elements(125);
      ct_core_CP_345_elements(124)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_345_elements(126);
      ct_core_CP_345_elements(115) <= phi_mux_reqs(1);
      phi_stmt_132_phi_seq_663 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_132_phi_seq_663") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_345_elements(110), 
          phi_sample_ack => ct_core_CP_345_elements(111), 
          phi_update_req => ct_core_CP_345_elements(112), 
          phi_update_ack => ct_core_CP_345_elements(113), 
          phi_mux_ack => ct_core_CP_345_elements(118), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_375_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ct_core_CP_345_elements(7);
        preds(1)  <= ct_core_CP_345_elements(8);
        entry_tmerge_375 : transition_merge -- 
          generic map(name => " entry_tmerge_375")
          port map (preds => preds, symbol_out => ct_core_CP_345_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_259_wire : std_logic_vector(15 downto 0);
    signal MUX_281_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_201_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_255_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_277_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_304_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_187_187_delayed_1_0_193 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_283_283_delayed_1_0_295 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_124 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_100 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_100_126_buffered : std_logic_vector(15 downto 0);
    signal add_dest_dim1_128 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_105 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_105_130_buffered : std_logic_vector(15 downto 0);
    signal add_out_161 : std_logic_vector(15 downto 0);
    signal add_src_132 : std_logic_vector(31 downto 0);
    signal add_src_init_109 : std_logic_vector(31 downto 0);
    signal cmp_dim0_204 : std_logic_vector(0 downto 0);
    signal cmp_dim1_198 : std_logic_vector(0 downto 0);
    signal cmp_dim2_188 : std_logic_vector(0 downto 0);
    signal continue_flag_306 : std_logic_vector(0 downto 0);
    signal dim0_end_300 : std_logic_vector(0 downto 0);
    signal dim2_limit_180 : std_logic_vector(15 downto 0);
    signal dim2_limit_180_delayed_1_0_183 : std_logic_vector(15 downto 0);
    signal done_175 : std_logic_vector(0 downto 0);
    signal i1_166 : std_logic_vector(63 downto 0);
    signal input_dim0_112 : std_logic_vector(15 downto 0);
    signal input_dim0_init_82 : std_logic_vector(15 downto 0);
    signal input_dim1_116 : std_logic_vector(15 downto 0);
    signal input_dim1_init_86 : std_logic_vector(15 downto 0);
    signal input_dim2_120 : std_logic_vector(15 downto 0);
    signal input_dim2_init_90 : std_logic_vector(15 downto 0);
    signal konst_159_wire_constant : std_logic_vector(15 downto 0);
    signal konst_178_wire_constant : std_logic_vector(15 downto 0);
    signal konst_191_wire_constant : std_logic_vector(15 downto 0);
    signal konst_207_wire_constant : std_logic_vector(15 downto 0);
    signal konst_212_wire_constant : std_logic_vector(15 downto 0);
    signal konst_222_wire_constant : std_logic_vector(15 downto 0);
    signal konst_250_wire_constant : std_logic_vector(31 downto 0);
    signal konst_272_wire_constant : std_logic_vector(15 downto 0);
    signal konst_279_wire_constant : std_logic_vector(15 downto 0);
    signal konst_293_wire_constant : std_logic_vector(15 downto 0);
    signal konst_93_wire_constant : std_logic_vector(15 downto 0);
    signal nao1_146 : std_logic_vector(15 downto 0);
    signal nao2_151 : std_logic_vector(15 downto 0);
    signal nao3_156 : std_logic_vector(15 downto 0);
    signal nao_141 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_268 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_268_127_buffered : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_262 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_262_131_buffered : std_logic_vector(15 downto 0);
    signal next_add_src_252 : std_logic_vector(31 downto 0);
    signal next_add_src_252_135_buffered : std_logic_vector(31 downto 0);
    signal next_input_dim0_290 : std_logic_vector(15 downto 0);
    signal next_input_dim0_290_115_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim1_284 : std_logic_vector(15 downto 0);
    signal next_input_dim1_284_119_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim2_274 : std_logic_vector(15 downto 0);
    signal next_input_dim2_274_123_buffered : std_logic_vector(15 downto 0);
    signal nid1_true1_229 : std_logic_vector(15 downto 0);
    signal nid1_true2_234 : std_logic_vector(15 downto 0);
    signal nid1_true3_233_delayed_1_0_242 : std_logic_vector(15 downto 0);
    signal nid1_true3_239 : std_logic_vector(15 downto 0);
    signal nid1_true4_247 : std_logic_vector(15 downto 0);
    signal nid1_true_224 : std_logic_vector(15 downto 0);
    signal nid2_false1_219 : std_logic_vector(15 downto 0);
    signal nid2_false_214 : std_logic_vector(15 downto 0);
    signal nid2_true_209 : std_logic_vector(15 downto 0);
    signal pad_95 : std_logic_vector(15 downto 0);
    signal type_cast_164_wire : std_logic_vector(31 downto 0);
    signal type_cast_169_169_delayed_15_0_170 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    add_src_init_109 <= "00000000000000000000000000000000";
    input_dim0_init_82 <= "0000000000000000";
    input_dim1_init_86 <= "0000000000000000";
    input_dim2_init_90 <= "0000000000000000";
    konst_159_wire_constant <= "0000000000000011";
    konst_178_wire_constant <= "0000000000001000";
    konst_191_wire_constant <= "0000000000000001";
    konst_207_wire_constant <= "0000000000001000";
    konst_212_wire_constant <= "0000000000000001";
    konst_222_wire_constant <= "0000000000000001";
    konst_250_wire_constant <= "00000000000000000000000000000001";
    konst_272_wire_constant <= "0000000000000000";
    konst_279_wire_constant <= "0000000000000000";
    konst_293_wire_constant <= "0000000000000001";
    konst_93_wire_constant <= "0000000000000001";
    phi_stmt_112: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim0_init_82 & next_input_dim0_290_115_buffered;
      req <= phi_stmt_112_req_0 & phi_stmt_112_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_112",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_112_ack_0,
          idata => idata,
          odata => input_dim0_112,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_112
    phi_stmt_116: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim1_init_86 & next_input_dim1_284_119_buffered;
      req <= phi_stmt_116_req_0 & phi_stmt_116_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_116",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_116_ack_0,
          idata => idata,
          odata => input_dim1_116,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_116
    phi_stmt_120: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim2_init_90 & next_input_dim2_274_123_buffered;
      req <= phi_stmt_120_req_0 & phi_stmt_120_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_120",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_120_ack_0,
          idata => idata,
          odata => input_dim2_120,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_120
    phi_stmt_124: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_dest_dim0_init_100_126_buffered & next_add_dest_dim0_268_127_buffered;
      req <= phi_stmt_124_req_0 & phi_stmt_124_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_124",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_124_ack_0,
          idata => idata,
          odata => add_dest_dim0_124,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_124
    phi_stmt_128: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_dest_dim1_init_105_130_buffered & next_add_dest_dim1_262_131_buffered;
      req <= phi_stmt_128_req_0 & phi_stmt_128_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_128",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_128_ack_0,
          idata => idata,
          odata => add_dest_dim1_128,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_128
    phi_stmt_132: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_src_init_109 & next_add_src_252_135_buffered;
      req <= phi_stmt_132_req_0 & phi_stmt_132_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_132",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_132_ack_0,
          idata => idata,
          odata => add_src_132,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_132
    -- flow-through select operator MUX_259_inst
    MUX_259_wire <= nid1_true4_247 when (cmp_dim1_198(0) /=  '0') else nid2_false1_219;
    -- flow-through select operator MUX_261_inst
    next_add_dest_dim1_262 <= MUX_259_wire when (NOT_u1_u1_255_wire(0) /=  '0') else add_dest_dim1_128;
    -- flow-through select operator MUX_267_inst
    next_add_dest_dim0_268 <= nid1_true1_229 when (cmp_dim0_204(0) /=  '0') else add_dest_dim0_124;
    -- flow-through select operator MUX_273_inst
    next_input_dim2_274 <= nid2_true_209 when (cmp_dim2_188(0) /=  '0') else konst_272_wire_constant;
    -- flow-through select operator MUX_281_inst
    MUX_281_wire <= konst_279_wire_constant when (cmp_dim1_198(0) /=  '0') else nid2_false_214;
    -- flow-through select operator MUX_283_inst
    next_input_dim1_284 <= MUX_281_wire when (NOT_u1_u1_277_wire(0) /=  '0') else input_dim1_116;
    -- flow-through select operator MUX_289_inst
    next_input_dim0_290 <= nid1_true_224 when (cmp_dim0_204(0) /=  '0') else input_dim0_112;
    W_dim2_limit_180_delayed_1_0_181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_dim2_limit_180_delayed_1_0_181_inst_req_0;
      W_dim2_limit_180_delayed_1_0_181_inst_ack_0<= wack(0);
      rreq(0) <= W_dim2_limit_180_delayed_1_0_181_inst_req_1;
      W_dim2_limit_180_delayed_1_0_181_inst_ack_1<= rack(0);
      W_dim2_limit_180_delayed_1_0_181_inst : InterlockBuffer generic map ( -- 
        name => "W_dim2_limit_180_delayed_1_0_181_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => dim2_limit_180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => dim2_limit_180_delayed_1_0_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_nid1_true3_233_delayed_1_0_240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_nid1_true3_233_delayed_1_0_240_inst_req_0;
      W_nid1_true3_233_delayed_1_0_240_inst_ack_0<= wack(0);
      rreq(0) <= W_nid1_true3_233_delayed_1_0_240_inst_req_1;
      W_nid1_true3_233_delayed_1_0_240_inst_ack_1<= rack(0);
      W_nid1_true3_233_delayed_1_0_240_inst : InterlockBuffer generic map ( -- 
        name => "W_nid1_true3_233_delayed_1_0_240_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nid1_true3_239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nid1_true3_233_delayed_1_0_242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim0_init_100_126_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim0_init_100_126_buf_req_0;
      add_dest_dim0_init_100_126_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim0_init_100_126_buf_req_1;
      add_dest_dim0_init_100_126_buf_ack_1<= rack(0);
      add_dest_dim0_init_100_126_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim0_init_100_126_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0_init_100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim0_init_100_126_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim1_init_105_130_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim1_init_105_130_buf_req_0;
      add_dest_dim1_init_105_130_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim1_init_105_130_buf_req_1;
      add_dest_dim1_init_105_130_buf_ack_1<= rack(0);
      add_dest_dim1_init_105_130_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim1_init_105_130_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1_init_105,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim1_init_105_130_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim0_268_127_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim0_268_127_buf_req_0;
      next_add_dest_dim0_268_127_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim0_268_127_buf_req_1;
      next_add_dest_dim0_268_127_buf_ack_1<= rack(0);
      next_add_dest_dim0_268_127_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim0_268_127_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim0_268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim0_268_127_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim1_262_131_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim1_262_131_buf_req_0;
      next_add_dest_dim1_262_131_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim1_262_131_buf_req_1;
      next_add_dest_dim1_262_131_buf_ack_1<= rack(0);
      next_add_dest_dim1_262_131_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim1_262_131_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim1_262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim1_262_131_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_src_252_135_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_src_252_135_buf_req_0;
      next_add_src_252_135_buf_ack_0<= wack(0);
      rreq(0) <= next_add_src_252_135_buf_req_1;
      next_add_src_252_135_buf_ack_1<= rack(0);
      next_add_src_252_135_buf : InterlockBuffer generic map ( -- 
        name => "next_add_src_252_135_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_src_252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_src_252_135_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim0_290_115_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim0_290_115_buf_req_0;
      next_input_dim0_290_115_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim0_290_115_buf_req_1;
      next_input_dim0_290_115_buf_ack_1<= rack(0);
      next_input_dim0_290_115_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim0_290_115_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim0_290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim0_290_115_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim1_284_119_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim1_284_119_buf_req_0;
      next_input_dim1_284_119_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim1_284_119_buf_req_1;
      next_input_dim1_284_119_buf_ack_1<= rack(0);
      next_input_dim1_284_119_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim1_284_119_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim1_284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim1_284_119_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim2_274_123_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim2_274_123_buf_req_0;
      next_input_dim2_274_123_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim2_274_123_buf_req_1;
      next_input_dim2_274_123_buf_ack_1<= rack(0);
      next_input_dim2_274_123_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim2_274_123_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim2_274,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim2_274_123_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_164_inst
    process(add_src_132) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_src_132(31 downto 0);
      type_cast_164_wire <= tmp_var; -- 
    end process;
    type_cast_169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_169_inst_req_0;
      type_cast_169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_169_inst_req_1;
      type_cast_169_inst_ack_1<= rack(0);
      type_cast_169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_169_inst",
        buffer_size => 15,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_out_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_169_169_delayed_15_0_170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_110_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_306;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_110_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_110_branch_req_0,
          ack0 => do_while_stmt_110_branch_ack_0,
          ack1 => do_while_stmt_110_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_145_inst
    process(nao_141, add_dest_dim1_128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nao_141, add_dest_dim1_128, tmp_var);
      nao1_146 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_155_inst
    process(input_dim2_120, nao2_151) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_120, nao2_151, tmp_var);
      nao3_156 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_208_inst
    process(input_dim2_120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_120, konst_207_wire_constant, tmp_var);
      nid2_true_209 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_213_inst
    process(input_dim1_116) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1_116, konst_212_wire_constant, tmp_var);
      nid2_false_214 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_218_inst
    process(add_dest_dim1_128, stride_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim1_128, stride_buffer, tmp_var);
      nid2_false1_219 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_223_inst
    process(input_dim0_112) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0_112, konst_222_wire_constant, tmp_var);
      nid1_true_224 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_228_inst
    process(add_dest_dim0_124, stride_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim0_124, stride_buffer, tmp_var);
      nid1_true1_229 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_94_inst
    process(padding_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(padding_buffer, konst_93_wire_constant, tmp_var);
      pad_95 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_251_inst
    process(add_src_132) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_src_132, konst_250_wire_constant, tmp_var);
      next_add_src_252 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_203_inst
    process(NOT_u1_u1_201_wire, cmp_dim1_198) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_201_wire, cmp_dim1_198, tmp_var);
      cmp_dim0_204 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_197_inst
    process(input_dim1_116, SUB_u16_u16_187_187_delayed_1_0_193) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1_116, SUB_u16_u16_187_187_delayed_1_0_193, tmp_var);
      cmp_dim1_198 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_160_inst
    process(nao3_156) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nao3_156, konst_159_wire_constant, tmp_var);
      add_out_161 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_140_inst
    process(out_d1_buffer, add_dest_dim0_124) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d1_buffer, add_dest_dim0_124, tmp_var);
      nao_141 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_150_inst
    process(out_d2_buffer, nao1_146) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d2_buffer, nao1_146, tmp_var);
      nao2_151 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_233_inst
    process(stride_buffer, inp_d1_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(stride_buffer, inp_d1_buffer, tmp_var);
      nid1_true2_234 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_201_inst
    process(cmp_dim2_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_188, tmp_var);
      NOT_u1_u1_201_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_255_inst
    process(cmp_dim2_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_188, tmp_var);
      NOT_u1_u1_255_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_277_inst
    process(cmp_dim2_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_188, tmp_var);
      NOT_u1_u1_277_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_304_inst
    process(cmp_dim0_204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim0_204, tmp_var);
      NOT_u1_u1_304_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_305_inst
    process(dim0_end_300, NOT_u1_u1_304_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(dim0_end_300, NOT_u1_u1_304_wire, tmp_var);
      continue_flag_306 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_104_inst
    process(ker_d2_buffer, pad_95) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(ker_d2_buffer, pad_95, tmp_var);
      add_dest_dim1_init_105 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_179_inst
    process(inp_d2_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(inp_d2_buffer, konst_178_wire_constant, tmp_var);
      dim2_limit_180 <= tmp_var; --
    end process;
    -- shared split operator group (22) : SUB_u16_u16_192_inst 
    ApIntSub_group_22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d1_buffer;
      SUB_u16_u16_187_187_delayed_1_0_193 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_192_inst_req_0;
      SUB_u16_u16_192_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_192_inst_req_1;
      SUB_u16_u16_192_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_22_gI: SplitGuardInterface generic map(name => "ApIntSub_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- binary operator SUB_u16_u16_238_inst
    process(nid1_true2_234, stride_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(nid1_true2_234, stride_buffer, tmp_var);
      nid1_true3_239 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_246_inst
    process(add_dest_dim1_128, nid1_true3_233_delayed_1_0_242) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add_dest_dim1_128, nid1_true3_233_delayed_1_0_242, tmp_var);
      nid1_true4_247 <= tmp_var; --
    end process;
    -- shared split operator group (25) : SUB_u16_u16_294_inst 
    ApIntSub_group_25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d0_buffer;
      SUB_u16_u16_283_283_delayed_1_0_295 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_294_inst_req_0;
      SUB_u16_u16_294_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_294_inst_req_1;
      SUB_u16_u16_294_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_25_gI: SplitGuardInterface generic map(name => "ApIntSub_group_25_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- binary operator SUB_u16_u16_99_inst
    process(ker_d1_buffer, pad_95) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(ker_d1_buffer, pad_95, tmp_var);
      add_dest_dim0_init_100 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_187_inst
    process(input_dim2_120, dim2_limit_180_delayed_1_0_183) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim2_120, dim2_limit_180_delayed_1_0_183, tmp_var);
      cmp_dim2_188 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_299_inst
    process(input_dim0_112, SUB_u16_u16_283_283_delayed_1_0_295) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim0_112, SUB_u16_u16_283_283_delayed_1_0_295, tmp_var);
      dim0_end_300 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_166_call 
    readModule1_call_group_0: Block -- 
      signal data_in: std_logic_vector(39 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 15);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_166_call_req_0;
      call_stmt_166_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_166_call_req_1;
      call_stmt_166_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      readModule1_call_group_0_gI: SplitGuardInterface generic map(name => "readModule1_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index1_buffer & type_cast_164_wire;
      i1_166 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 40,
        owidth => 40,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => readModule1_call_reqs(0),
          ackR => readModule1_call_acks(0),
          dataR => readModule1_call_data(39 downto 0),
          tagR => readModule1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => readModule1_return_acks(0), -- cross-over
          ackL => readModule1_return_reqs(0), -- cross-over
          dataL => readModule1_return_data(63 downto 0),
          tagL => readModule1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_175_call 
    writeModule1_call_group_1: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 9);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_175_call_req_0;
      call_stmt_175_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_175_call_req_1;
      call_stmt_175_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeModule1_call_group_1_gI: SplitGuardInterface generic map(name => "writeModule1_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index3_buffer & type_cast_169_169_delayed_15_0_170 & i1_166;
      done_175 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeModule1_call_reqs(0),
          ackR => writeModule1_call_acks(0),
          dataR => writeModule1_call_data(103 downto 0),
          tagR => writeModule1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeModule1_return_acks(0), -- cross-over
          ackL => writeModule1_return_reqs(0), -- cross-over
          dataL => writeModule1_return_data(0 downto 0),
          tagL => writeModule1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end ct_core_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readModule1;
architecture readModule1_arch of readModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 40)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  -- output port buffer signals
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  signal readModule1_CP_34_start: Boolean;
  signal readModule1_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_32_index_0_scale_req_0 : boolean;
  signal ptr_deref_37_load_0_req_0 : boolean;
  signal array_obj_ref_32_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_32_index_0_scale_req_1 : boolean;
  signal array_obj_ref_32_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_32_index_sum_1_req_0 : boolean;
  signal array_obj_ref_32_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_32_index_sum_1_req_1 : boolean;
  signal array_obj_ref_32_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_32_index_offset_req_0 : boolean;
  signal array_obj_ref_32_index_offset_ack_0 : boolean;
  signal array_obj_ref_32_index_offset_req_1 : boolean;
  signal array_obj_ref_32_index_offset_ack_1 : boolean;
  signal addr_of_33_final_reg_req_0 : boolean;
  signal addr_of_33_final_reg_ack_0 : boolean;
  signal addr_of_33_final_reg_req_1 : boolean;
  signal addr_of_33_final_reg_ack_1 : boolean;
  signal ptr_deref_37_load_0_ack_0 : boolean;
  signal ptr_deref_37_load_0_req_1 : boolean;
  signal ptr_deref_37_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readModule1_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 40) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(tag_length + 39 downto 40) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 39 downto 40);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 3) := (0 => 8,1 => 8,2 => 1,3 => 8);
    constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 8);
    constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 4); -- 
  begin -- 
    preds <= index_update_enable & address_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readModule1_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readModule1_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= data_buffer;
  data <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  data_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "data_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_data_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => data_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readModule1_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readModule1_CP_34: Block -- control-path 
    signal readModule1_CP_34_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    readModule1_CP_34_elements(0) <= readModule1_CP_34_start;
    readModule1_CP_34_symbol <= readModule1_CP_34_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	17 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resized_0
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_computed_0
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resized_2
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scaled_2
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_computed_2
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/$exit
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/index_resize_req
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/$exit
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/scale_rename_ack
      -- 
    readModule1_CP_34_elements(1) <= readModule1_CP_34_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	27 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_34_to_assign_stmt_38/index_update_enable
      -- CP-element group 2: 	 assign_stmt_34_to_assign_stmt_38/index_update_enable_out
      -- 
    readModule1_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readModule1_CP_34_elements(8);
      gj_readModule1_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	28 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_34_to_assign_stmt_38/address_update_enable
      -- CP-element group 3: 	 assign_stmt_34_to_assign_stmt_38/address_update_enable_out
      -- 
    readModule1_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readModule1_CP_34_elements(15);
      gj_readModule1_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	29 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	23 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_34_to_assign_stmt_38/data_update_enable
      -- CP-element group 4: 	 assign_stmt_34_to_assign_stmt_38/data_update_enable_in
      -- 
    readModule1_CP_34_elements(4) <= readModule1_CP_34_elements(29);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	20 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_sample_start_
      -- CP-element group 5: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/$entry
      -- CP-element group 5: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/req
      -- 
    req_121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(5), ack => addr_of_33_final_reg_req_0); -- 
    readModule1_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(7) & readModule1_CP_34_elements(20);
      gj_readModule1_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	24 
    -- CP-element group 6: 	21 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_update_start_
      -- CP-element group 6: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/$entry
      -- CP-element group 6: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/req
      -- 
    req_126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(6), ack => addr_of_33_final_reg_req_1); -- 
    readModule1_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(24) & readModule1_CP_34_elements(21);
      gj_readModule1_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	16 
    -- CP-element group 7: 	19 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	17 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_root_address_calculated
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_offset_calculated
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/$entry
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/$exit
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/sum_rename_req
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/sum_rename_ack
      -- 
    readModule1_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(16) & readModule1_CP_34_elements(19);
      gj_readModule1_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	15 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scaled_0
      -- 
    readModule1_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(12) & readModule1_CP_34_elements(15);
      gj_readModule1_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/rr
      -- CP-element group 9: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_sample_start
      -- 
    rr_67_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_67_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(9), ack => array_obj_ref_32_index_0_scale_req_0); -- 
    readModule1_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(11);
      gj_readModule1_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_update_start
      -- CP-element group 10: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/$entry
      -- CP-element group 10: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/cr
      -- 
    cr_72_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_72_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(10), ack => array_obj_ref_32_index_0_scale_req_1); -- 
    readModule1_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(12);
      gj_readModule1_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	26 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_sample_complete
      -- CP-element group 11: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/ra
      -- 
    ra_68_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_0_scale_ack_0, ack => readModule1_CP_34_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_update_complete
      -- CP-element group 12: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/$exit
      -- CP-element group 12: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/ca
      -- 
    ca_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_0_scale_ack_1, ack => readModule1_CP_34_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: 	1 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_sample_start
      -- CP-element group 13: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/rr
      -- 
    rr_94_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_94_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(13), ack => array_obj_ref_32_index_sum_1_req_0); -- 
    readModule1_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 8,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(8) & readModule1_CP_34_elements(1) & readModule1_CP_34_elements(15);
      gj_readModule1_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_update_start
      -- CP-element group 14: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/$entry
      -- CP-element group 14: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/cr
      -- 
    cr_99_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_99_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(14), ack => array_obj_ref_32_index_sum_1_req_1); -- 
    readModule1_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(16) & readModule1_CP_34_elements(18);
      gj_readModule1_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	26 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	8 
    -- CP-element group 15: 	13 
    -- CP-element group 15: 	3 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_sample_complete
      -- CP-element group 15: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/ra
      -- 
    ra_95_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_sum_1_ack_0, ack => readModule1_CP_34_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: 	18 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_update_complete
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/$exit
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/ca
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/$entry
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/req
      -- 
    ca_100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_sum_1_ack_1, ack => readModule1_CP_34_elements(16)); -- 
    req_106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(16), ack => array_obj_ref_32_index_offset_req_0); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	7 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_update_start
      -- CP-element group 17: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/req
      -- 
    req_111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(17), ack => array_obj_ref_32_index_offset_req_1); -- 
    readModule1_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(7) & readModule1_CP_34_elements(20);
      gj_readModule1_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	26 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/ack
      -- 
    ack_107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_offset_ack_0, ack => readModule1_CP_34_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	7 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/ack
      -- 
    ack_112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_offset_ack_1, ack => readModule1_CP_34_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	5 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	5 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_sample_completed_
      -- CP-element group 20: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/$exit
      -- CP-element group 20: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/ack
      -- 
    ack_122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_33_final_reg_ack_0, ack => readModule1_CP_34_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	6 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_update_completed_
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/ack
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_address_resized
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/root_register_ack
      -- 
    ack_127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_33_final_reg_ack_1, ack => readModule1_CP_34_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/$entry
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/$entry
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/rr
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_sample_start_
      -- 
    rr_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(22), ack => ptr_deref_37_load_0_req_0); -- 
    readModule1_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(21) & readModule1_CP_34_elements(24);
      gj_readModule1_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	4 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_update_start_
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/$entry
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/$entry
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/$entry
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/cr
      -- 
    cr_171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(23), ack => ptr_deref_37_load_0_req_1); -- 
    readModule1_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(4) & readModule1_CP_34_elements(25);
      gj_readModule1_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	6 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/$exit
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_sample_completed_
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/ra
      -- 
    ra_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_37_load_0_ack_0, ack => readModule1_CP_34_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_update_completed_
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/$entry
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/merge_req
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/merge_ack
      -- 
    ca_172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_37_load_0_ack_1, ack => readModule1_CP_34_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	11 
    -- CP-element group 26: 	25 
    -- CP-element group 26: 	15 
    -- CP-element group 26: 	18 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	30 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 assign_stmt_34_to_assign_stmt_38/$exit
      -- 
    readModule1_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 8,1 => 8,2 => 8,3 => 8);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(11) & readModule1_CP_34_elements(25) & readModule1_CP_34_elements(15) & readModule1_CP_34_elements(18);
      gj_readModule1_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  place  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 index_update_enable
      -- 
    readModule1_CP_34_elements(27) <= readModule1_CP_34_elements(2);
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	3 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 address_update_enable
      -- 
    readModule1_CP_34_elements(28) <= readModule1_CP_34_elements(3);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	4 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 data_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	26 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    readModule1_CP_34_elements(30) <= readModule1_CP_34_elements(26);
    --  hookup: inputs to control-path 
    readModule1_CP_34_elements(29) <= data_update_enable;
    -- hookup: output from control-path 
    index_update_enable <= readModule1_CP_34_elements(27);
    address_update_enable <= readModule1_CP_34_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_address_31_resized : std_logic_vector(15 downto 0);
    signal R_address_31_scaled : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_index_partial_sum_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_root_address : std_logic_vector(15 downto 0);
    signal ptr_34 : std_logic_vector(31 downto 0);
    signal ptr_deref_37_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_37_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_37_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_37_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_37_word_offset_0 : std_logic_vector(15 downto 0);
    signal type_cast_28_resized : std_logic_vector(15 downto 0);
    signal type_cast_28_scaled : std_logic_vector(15 downto 0);
    signal type_cast_28_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_32_constant_part_of_offset <= "0000000000000000";
    array_obj_ref_32_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_32_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_32_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_32_resized_base_address <= "0000000000000000";
    ptr_deref_37_word_offset_0 <= "0000000000000000";
    addr_of_33_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_33_final_reg_req_0;
      addr_of_33_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_33_final_reg_req_1;
      addr_of_33_final_reg_ack_1<= rack(0);
      addr_of_33_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_33_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_32_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_34,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_28_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := index_buffer(7 downto 0);
      type_cast_28_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_32_index_0_resize
    process(type_cast_28_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_28_wire;
      ov := iv(15 downto 0);
      type_cast_28_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_32_index_2_rename
    process(R_address_31_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_31_resized;
      ov(15 downto 0) := iv;
      R_address_31_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_32_index_2_resize
    process(address_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_buffer;
      ov := iv(15 downto 0);
      R_address_31_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_32_root_address_inst
    process(array_obj_ref_32_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_32_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_32_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_addr_0
    process(ptr_deref_37_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_37_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_37_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_base_resize
    process(ptr_34) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_34;
      ov := iv(15 downto 0);
      ptr_deref_37_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_gather_scatter
    process(ptr_deref_37_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_37_data_0;
      ov(63 downto 0) := iv;
      data_buffer <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_root_address_inst
    process(ptr_deref_37_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_37_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_37_root_address <= ov(15 downto 0);
      --
    end process;
    -- shared split operator group (0) : array_obj_ref_32_index_0_scale 
    ApIntMul_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_28_resized;
      type_cast_28_scaled <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_32_index_0_scale_req_0;
      array_obj_ref_32_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_32_index_0_scale_req_1;
      array_obj_ref_32_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_0_gI: SplitGuardInterface generic map(name => "ApIntMul_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0100000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_32_index_offset 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_32_index_partial_sum_1;
      array_obj_ref_32_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_32_index_offset_req_0;
      array_obj_ref_32_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_32_index_offset_req_1;
      array_obj_ref_32_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_32_index_sum_1 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_31_scaled & type_cast_28_scaled;
      array_obj_ref_32_index_partial_sum_1 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_32_index_sum_1_req_0;
      array_obj_ref_32_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_32_index_sum_1_req_1;
      array_obj_ref_32_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared load operator group (0) : ptr_deref_37_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_37_load_0_req_0;
      ptr_deref_37_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_37_load_0_req_1;
      ptr_deref_37_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_37_word_address_0;
      ptr_deref_37_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(15 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end readModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_13_inst_req_0 : boolean;
  signal WPIPE_timer_req_13_inst_ack_0 : boolean;
  signal WPIPE_timer_req_13_inst_req_1 : boolean;
  signal WPIPE_timer_req_13_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_18_inst_req_0 : boolean;
  signal RPIPE_timer_resp_18_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_18_inst_req_1 : boolean;
  signal RPIPE_timer_resp_18_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/$entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_sample_start_
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/req
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_18_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_13_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_sample_completed_
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_update_start_
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/ack
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/$entry
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_13_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_13_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_update_completed_
      -- CP-element group 2: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/$exit
      -- CP-element group 2: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_13_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_sample_completed_
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_update_start_
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/ra
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/$entry
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_18_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_18_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_update_completed_
      -- CP-element group 4: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/$exit
      -- CP-element group 4: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_18_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_16_to_assign_stmt_19/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(2) & timer_CP_0_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_15_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_15_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_18_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_18_inst_req_0;
      RPIPE_timer_resp_18_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_18_inst_req_1;
      RPIPE_timer_resp_18_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_13_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_13_inst_req_0;
      WPIPE_timer_req_13_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_13_inst_req_1;
      WPIPE_timer_req_13_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_15_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_3687_start: Boolean;
  signal timerDaemon_CP_3687_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1580_branch_req_0 : boolean;
  signal phi_stmt_1582_req_1 : boolean;
  signal phi_stmt_1582_req_0 : boolean;
  signal phi_stmt_1582_ack_0 : boolean;
  signal nCOUNTER_1595_1586_buf_req_0 : boolean;
  signal nCOUNTER_1595_1586_buf_ack_0 : boolean;
  signal nCOUNTER_1595_1586_buf_req_1 : boolean;
  signal nCOUNTER_1595_1586_buf_ack_1 : boolean;
  signal RPIPE_timer_req_1589_inst_req_0 : boolean;
  signal RPIPE_timer_req_1589_inst_ack_0 : boolean;
  signal RPIPE_timer_req_1589_inst_req_1 : boolean;
  signal RPIPE_timer_req_1589_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_1597_inst_req_0 : boolean;
  signal WPIPE_timer_resp_1597_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_1597_inst_req_1 : boolean;
  signal WPIPE_timer_resp_1597_inst_ack_1 : boolean;
  signal do_while_stmt_1580_branch_ack_0 : boolean;
  signal do_while_stmt_1580_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_3687_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3687_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_3687_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3687_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_3687: Block -- control-path 
    signal timerDaemon_CP_3687_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_3687_elements(0) <= timerDaemon_CP_3687_start;
    timerDaemon_CP_3687_symbol <= timerDaemon_CP_3687_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1579/$entry
      -- CP-element group 0: 	 branch_block_stmt_1579/branch_block_stmt_1579__entry__
      -- CP-element group 0: 	 branch_block_stmt_1579/do_while_stmt_1580__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1579/$exit
      -- CP-element group 1: 	 branch_block_stmt_1579/branch_block_stmt_1579__exit__
      -- CP-element group 1: 	 branch_block_stmt_1579/do_while_stmt_1580__exit__
      -- 
    timerDaemon_CP_3687_elements(1) <= timerDaemon_CP_3687_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1579/do_while_stmt_1580/$entry
      -- CP-element group 2: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580__entry__
      -- 
    timerDaemon_CP_3687_elements(2) <= timerDaemon_CP_3687_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580__exit__
      -- 
    -- Element group timerDaemon_CP_3687_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_back
      -- 
    -- Element group timerDaemon_CP_3687_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1579/do_while_stmt_1580/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_taken/$entry
      -- 
    timerDaemon_CP_3687_elements(5) <= timerDaemon_CP_3687_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_body_done
      -- 
    timerDaemon_CP_3687_elements(6) <= timerDaemon_CP_3687_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_3687_elements(7) <= timerDaemon_CP_3687_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_3687_elements(8) <= timerDaemon_CP_3687_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1587_sample_start_
      -- 
    -- Element group timerDaemon_CP_3687_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/condition_evaluated
      -- 
    condition_evaluated_3711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(10), ack => do_while_stmt_1580_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(40) & timerDaemon_CP_3687_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(9) & timerDaemon_CP_3687_elements(15) & timerDaemon_CP_3687_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1587_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(35) & timerDaemon_CP_3687_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(32) & timerDaemon_CP_3687_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(36) & timerDaemon_CP_3687_elements(18);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(9) & timerDaemon_CP_3687_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(9) & timerDaemon_CP_3687_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_3687_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	37 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_3687_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_loopback_trigger
      -- 
    timerDaemon_CP_3687_elements(19) <= timerDaemon_CP_3687_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_loopback_sample_req_ps
      -- 
    phi_stmt_1582_loopback_sample_req_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1582_loopback_sample_req_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(20), ack => phi_stmt_1582_req_1); -- 
    -- Element group timerDaemon_CP_3687_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_entry_trigger
      -- 
    timerDaemon_CP_3687_elements(21) <= timerDaemon_CP_3687_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_entry_sample_req_ps
      -- 
    phi_stmt_1582_entry_sample_req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1582_entry_sample_req_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(22), ack => phi_stmt_1582_req_0); -- 
    -- Element group timerDaemon_CP_3687_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1582_phi_mux_ack_ps
      -- 
    phi_stmt_1582_phi_mux_ack_3732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1582_ack_0, ack => timerDaemon_CP_3687_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_sample_completed_
      -- 
    -- Element group timerDaemon_CP_3687_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_update_start_
      -- 
    -- Element group timerDaemon_CP_3687_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_update_completed__ps
      -- 
    timerDaemon_CP_3687_elements(26) <= timerDaemon_CP_3687_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/type_cast_1585_update_completed_
      -- 
    -- Element group timerDaemon_CP_3687_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_3687_elements(25), ack => timerDaemon_CP_3687_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Sample/req
      -- 
    req_3753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(28), ack => nCOUNTER_1595_1586_buf_req_0); -- 
    -- Element group timerDaemon_CP_3687_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Update/req
      -- 
    req_3758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(29), ack => nCOUNTER_1595_1586_buf_req_1); -- 
    -- Element group timerDaemon_CP_3687_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Sample/ack
      -- 
    ack_3754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1595_1586_buf_ack_0, ack => timerDaemon_CP_3687_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/R_nCOUNTER_1586_Update/ack
      -- 
    ack_3759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1595_1586_buf_ack_1, ack => timerDaemon_CP_3687_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1587_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(9) & timerDaemon_CP_3687_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Sample/rr
      -- 
    rr_3772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(33), ack => RPIPE_timer_req_1589_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(11) & timerDaemon_CP_3687_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Update/cr
      -- 
    cr_3777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(34), ack => RPIPE_timer_req_1589_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(35) & timerDaemon_CP_3687_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Sample/ra
      -- 
    ra_3773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1589_inst_ack_0, ack => timerDaemon_CP_3687_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/phi_stmt_1587_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/RPIPE_timer_req_1589_Update/ca
      -- 
    ca_3778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1589_inst_ack_1, ack => timerDaemon_CP_3687_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Sample/req
      -- 
    req_3786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(37), ack => WPIPE_timer_resp_1597_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(36) & timerDaemon_CP_3687_elements(18) & timerDaemon_CP_3687_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Update/req
      -- 
    ack_3787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1597_inst_ack_0, ack => timerDaemon_CP_3687_elements(38)); -- 
    req_3791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3687_elements(38), ack => WPIPE_timer_resp_1597_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/WPIPE_timer_resp_1597_Update/ack
      -- 
    ack_3792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1597_inst_ack_1, ack => timerDaemon_CP_3687_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_3687_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_3687_elements(9), ack => timerDaemon_CP_3687_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1579/do_while_stmt_1580/do_while_stmt_1580_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3687_elements(39) & timerDaemon_CP_3687_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3687_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_exit/ack
      -- 
    ack_3797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1580_branch_ack_0, ack => timerDaemon_CP_3687_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1579/do_while_stmt_1580/loop_taken/ack
      -- 
    ack_3801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1580_branch_ack_1, ack => timerDaemon_CP_3687_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1579/do_while_stmt_1580/$exit
      -- 
    timerDaemon_CP_3687_elements(44) <= timerDaemon_CP_3687_elements(3);
    timerDaemon_do_while_stmt_1580_terminator_3802: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1580_terminator_3802", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_3687_elements(6),loop_continue => timerDaemon_CP_3687_elements(43),loop_terminate => timerDaemon_CP_3687_elements(42),loop_back => timerDaemon_CP_3687_elements(4),loop_exit => timerDaemon_CP_3687_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1582_phi_seq_3760_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_3687_elements(21);
      timerDaemon_CP_3687_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_3687_elements(24);
      timerDaemon_CP_3687_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_3687_elements(26);
      timerDaemon_CP_3687_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_3687_elements(19);
      timerDaemon_CP_3687_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_3687_elements(30);
      timerDaemon_CP_3687_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_3687_elements(31);
      timerDaemon_CP_3687_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1582_phi_seq_3760 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1582_phi_seq_3760") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_3687_elements(11), 
          phi_sample_ack => timerDaemon_CP_3687_elements(17), 
          phi_update_req => timerDaemon_CP_3687_elements(13), 
          phi_update_ack => timerDaemon_CP_3687_elements(18), 
          phi_mux_ack => timerDaemon_CP_3687_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3712_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_3687_elements(7);
        preds(1)  <= timerDaemon_CP_3687_elements(8);
        entry_tmerge_3712 : transition_merge -- 
          generic map(name => " entry_tmerge_3712")
          port map (preds => preds, symbol_out => timerDaemon_CP_3687_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1582 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1589_wire : std_logic_vector(0 downto 0);
    signal konst_1593_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1601_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1595 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1595_1586_buffered : std_logic_vector(63 downto 0);
    signal req_1587 : std_logic_vector(0 downto 0);
    signal type_cast_1585_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1593_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1601_wire_constant <= "1";
    type_cast_1585_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1582: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1585_wire_constant & nCOUNTER_1595_1586_buffered;
      req <= phi_stmt_1582_req_0 & phi_stmt_1582_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1582",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1582_ack_0,
          idata => idata,
          odata => COUNTER_1582,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1582
    nCOUNTER_1595_1586_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1595_1586_buf_req_0;
      nCOUNTER_1595_1586_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1595_1586_buf_req_1;
      nCOUNTER_1595_1586_buf_ack_1<= rack(0);
      nCOUNTER_1595_1586_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1595_1586_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1595_1586_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1587
    process(RPIPE_timer_req_1589_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1589_wire(0 downto 0);
      req_1587 <= tmp_var; -- 
    end process;
    do_while_stmt_1580_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1601_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1580_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1580_branch_req_0,
          ack0 => do_while_stmt_1580_branch_ack_0,
          ack1 => do_while_stmt_1580_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1594_inst
    process(COUNTER_1582) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1582, konst_1593_wire_constant, tmp_var);
      nCOUNTER_1595 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1589_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1589_inst_req_0;
      RPIPE_timer_req_1589_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1589_inst_req_1;
      RPIPE_timer_req_1589_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1589_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1597_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1597_inst_req_0;
      WPIPE_timer_resp_1597_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1597_inst_req_1;
      WPIPE_timer_resp_1597_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1587(0);
      data_in <= COUNTER_1582;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity writeModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : in  std_logic_vector(63 downto 0);
    done : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeModule1;
architecture writeModule1_arch of writeModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 104)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  -- output port buffer signals
  signal done_buffer :  std_logic_vector(0 downto 0);
  signal done_update_enable: Boolean;
  signal writeModule1_CP_181_start: Boolean;
  signal writeModule1_CP_181_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_51_index_0_scale_req_0 : boolean;
  signal array_obj_ref_51_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_51_index_0_scale_req_1 : boolean;
  signal array_obj_ref_51_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_51_index_sum_1_req_0 : boolean;
  signal array_obj_ref_51_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_51_index_sum_1_req_1 : boolean;
  signal array_obj_ref_51_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_51_index_offset_req_0 : boolean;
  signal array_obj_ref_51_index_offset_ack_0 : boolean;
  signal array_obj_ref_51_index_offset_req_1 : boolean;
  signal array_obj_ref_51_index_offset_ack_1 : boolean;
  signal addr_of_52_final_reg_req_0 : boolean;
  signal addr_of_52_final_reg_ack_0 : boolean;
  signal addr_of_52_final_reg_req_1 : boolean;
  signal addr_of_52_final_reg_ack_1 : boolean;
  signal ptr_deref_55_store_0_req_0 : boolean;
  signal ptr_deref_55_store_0_ack_0 : boolean;
  signal ptr_deref_55_store_0_req_1 : boolean;
  signal ptr_deref_55_store_0_ack_1 : boolean;
  signal BITSEL_u8_u1_61_inst_req_0 : boolean;
  signal BITSEL_u8_u1_61_inst_ack_0 : boolean;
  signal BITSEL_u8_u1_61_inst_req_1 : boolean;
  signal BITSEL_u8_u1_61_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeModule1_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 104) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(103 downto 40) <= data;
  data_buffer <= in_buffer_data_out(103 downto 40);
  in_buffer_data_in(tag_length + 103 downto 104) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 103 downto 104);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 8,1 => 8,2 => 8,3 => 1,4 => 8);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 8);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= index_update_enable & address_update_enable & data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeModule1_CP_181_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeModule1_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= done_buffer;
  done <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_181_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  done_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "done_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_done_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => done_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeModule1_CP_181_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_181_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeModule1_CP_181: Block -- control-path 
    signal writeModule1_CP_181_elements: BooleanArray(36 downto 0);
    -- 
  begin -- 
    writeModule1_CP_181_elements(0) <= writeModule1_CP_181_start;
    writeModule1_CP_181_symbol <= writeModule1_CP_181_elements(36);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	27 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	15 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resized_0
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_computed_0
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resized_2
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scaled_2
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_computed_2
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/$exit
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/index_resize_req
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/$exit
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/scale_rename_ack
      -- 
    writeModule1_CP_181_elements(1) <= writeModule1_CP_181_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	32 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_53_to_assign_stmt_62/index_update_enable
      -- CP-element group 2: 	 assign_stmt_53_to_assign_stmt_62/index_update_enable_out
      -- 
    writeModule1_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(29) & writeModule1_CP_181_elements(9);
      gj_writeModule1_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	16 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	33 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_53_to_assign_stmt_62/address_update_enable
      -- CP-element group 3: 	 assign_stmt_53_to_assign_stmt_62/address_update_enable_out
      -- 
    writeModule1_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_181_elements(16);
      gj_writeModule1_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	25 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	34 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_53_to_assign_stmt_62/data_update_enable
      -- CP-element group 4: 	 assign_stmt_53_to_assign_stmt_62/data_update_enable_out
      -- 
    writeModule1_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_181_elements(25);
      gj_writeModule1_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	35 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	28 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_53_to_assign_stmt_62/done_update_enable
      -- CP-element group 5: 	 assign_stmt_53_to_assign_stmt_62/done_update_enable_in
      -- 
    writeModule1_CP_181_elements(5) <= writeModule1_CP_181_elements(35);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	21 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_sample_start_
      -- CP-element group 6: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/$entry
      -- CP-element group 6: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/req
      -- 
    req_270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(6), ack => addr_of_52_final_reg_req_0); -- 
    writeModule1_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(8) & writeModule1_CP_181_elements(21);
      gj_writeModule1_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	25 
    -- CP-element group 7: 	22 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	22 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_update_start_
      -- CP-element group 7: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/$entry
      -- CP-element group 7: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/req
      -- 
    req_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(7), ack => addr_of_52_final_reg_req_1); -- 
    writeModule1_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(25) & writeModule1_CP_181_elements(22);
      gj_writeModule1_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	20 
    -- CP-element group 8: 	17 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_root_address_calculated
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_offset_calculated
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/$entry
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/$exit
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/sum_rename_ack
      -- 
    writeModule1_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 8);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(20) & writeModule1_CP_181_elements(17);
      gj_writeModule1_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	13 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	2 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scaled_0
      -- 
    writeModule1_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(13) & writeModule1_CP_181_elements(16);
      gj_writeModule1_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_sample_start
      -- CP-element group 10: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/rr
      -- 
    rr_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(10), ack => array_obj_ref_51_index_0_scale_req_0); -- 
    writeModule1_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(12);
      gj_writeModule1_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_update_start
      -- CP-element group 11: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/$entry
      -- CP-element group 11: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/cr
      -- 
    cr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(11), ack => array_obj_ref_51_index_0_scale_req_1); -- 
    writeModule1_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(13);
      gj_writeModule1_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_sample_complete
      -- CP-element group 12: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/ra
      -- 
    ra_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_0_scale_ack_0, ack => writeModule1_CP_181_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_update_complete
      -- CP-element group 13: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/$exit
      -- CP-element group 13: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/ca
      -- 
    ca_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_0_scale_ack_1, ack => writeModule1_CP_181_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_sample_start
      -- CP-element group 14: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/rr
      -- 
    rr_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(14), ack => array_obj_ref_51_index_sum_1_req_0); -- 
    writeModule1_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(9) & writeModule1_CP_181_elements(16);
      gj_writeModule1_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	1 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_update_start
      -- CP-element group 15: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/$entry
      -- CP-element group 15: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/cr
      -- 
    cr_248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(15), ack => array_obj_ref_51_index_sum_1_req_1); -- 
    writeModule1_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(17) & writeModule1_CP_181_elements(19);
      gj_writeModule1_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_sample_complete
      -- CP-element group 16: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/ra
      -- 
    ra_244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_sum_1_ack_0, ack => writeModule1_CP_181_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	8 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_update_complete
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/$exit
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/ca
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/req
      -- 
    ca_249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_sum_1_ack_1, ack => writeModule1_CP_181_elements(17)); -- 
    req_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(17), ack => array_obj_ref_51_index_offset_req_0); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_update_start
      -- CP-element group 18: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/$entry
      -- CP-element group 18: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/req
      -- 
    req_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(18), ack => array_obj_ref_51_index_offset_req_1); -- 
    writeModule1_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(8) & writeModule1_CP_181_elements(21);
      gj_writeModule1_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	31 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_sample_complete
      -- CP-element group 19: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/ack
      -- 
    ack_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_offset_ack_0, ack => writeModule1_CP_181_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	8 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/$exit
      -- CP-element group 20: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/ack
      -- 
    ack_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_offset_ack_1, ack => writeModule1_CP_181_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	6 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_sample_completed_
      -- CP-element group 21: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/$exit
      -- CP-element group 21: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/ack
      -- 
    ack_271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_52_final_reg_ack_0, ack => writeModule1_CP_181_elements(21)); -- 
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	7 
    -- CP-element group 22:  members (19) 
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_update_completed_
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/ack
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_address_calculated
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_address_calculated
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_root_address_calculated
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_address_resized
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/$entry
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/base_resize_req
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/base_resize_ack
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/$entry
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/sum_rename_req
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/sum_rename_ack
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/$entry
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/root_register_req
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/root_register_ack
      -- 
    ack_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_52_final_reg_ack_1, ack => writeModule1_CP_181_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: 	22 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_sample_start_
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/$exit
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/split_req
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/split_ack
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/rr
      -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(23), ack => ptr_deref_55_store_0_req_0); -- 
    writeModule1_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(22) & writeModule1_CP_181_elements(25);
      gj_writeModule1_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_update_start_
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/$entry
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/$entry
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/$entry
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/cr
      -- 
    cr_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(24), ack => ptr_deref_55_store_0_req_1); -- 
    writeModule1_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_181_elements(26);
      gj_writeModule1_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: 	7 
    -- CP-element group 25: 	4 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_sample_completed_
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/$exit
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/ra
      -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_55_store_0_ack_0, ack => writeModule1_CP_181_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_update_completed_
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/$exit
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/$exit
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/ca
      -- 
    ca_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_55_store_0_ack_1, ack => writeModule1_CP_181_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	1 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_sample_start_
      -- CP-element group 27: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/rr
      -- 
    rr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(27), ack => BITSEL_u8_u1_61_inst_req_0); -- 
    writeModule1_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(29);
      gj_writeModule1_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	5 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_update_start_
      -- CP-element group 28: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/$entry
      -- CP-element group 28: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/cr
      -- 
    cr_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(28), ack => BITSEL_u8_u1_61_inst_req_1); -- 
    writeModule1_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(5) & writeModule1_CP_181_elements(30);
      gj_writeModule1_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_sample_completed_
      -- CP-element group 29: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/$exit
      -- CP-element group 29: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/ra
      -- 
    ra_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_61_inst_ack_0, ack => writeModule1_CP_181_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_update_completed_
      -- CP-element group 30: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/$exit
      -- CP-element group 30: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/ca
      -- 
    ca_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_61_inst_ack_1, ack => writeModule1_CP_181_elements(30)); -- 
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	19 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	12 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 assign_stmt_53_to_assign_stmt_62/$exit
      -- 
    writeModule1_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 8,1 => 8,2 => 8,3 => 8,4 => 8);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(19) & writeModule1_CP_181_elements(16) & writeModule1_CP_181_elements(26) & writeModule1_CP_181_elements(12) & writeModule1_CP_181_elements(30);
      gj_writeModule1_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  place  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 index_update_enable
      -- 
    writeModule1_CP_181_elements(32) <= writeModule1_CP_181_elements(2);
    -- CP-element group 33:  place  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	3 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 address_update_enable
      -- 
    writeModule1_CP_181_elements(33) <= writeModule1_CP_181_elements(3);
    -- CP-element group 34:  place  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	4 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 data_update_enable
      -- 
    writeModule1_CP_181_elements(34) <= writeModule1_CP_181_elements(4);
    -- CP-element group 35:  place  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	5 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 done_update_enable
      -- 
    -- CP-element group 36:  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 $exit
      -- 
    writeModule1_CP_181_elements(36) <= writeModule1_CP_181_elements(31);
    --  hookup: inputs to control-path 
    writeModule1_CP_181_elements(35) <= done_update_enable;
    -- hookup: output from control-path 
    index_update_enable <= writeModule1_CP_181_elements(32);
    address_update_enable <= writeModule1_CP_181_elements(33);
    data_update_enable <= writeModule1_CP_181_elements(34);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_address_50_resized : std_logic_vector(15 downto 0);
    signal R_address_50_scaled : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_index_partial_sum_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_root_address : std_logic_vector(15 downto 0);
    signal konst_60_wire_constant : std_logic_vector(7 downto 0);
    signal ptr_53 : std_logic_vector(31 downto 0);
    signal ptr_deref_55_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_55_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_55_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_55_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_55_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_55_word_offset_0 : std_logic_vector(15 downto 0);
    signal type_cast_47_resized : std_logic_vector(15 downto 0);
    signal type_cast_47_scaled : std_logic_vector(15 downto 0);
    signal type_cast_47_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_51_constant_part_of_offset <= "0000000000000000";
    array_obj_ref_51_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_51_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_51_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_51_resized_base_address <= "0000000000000000";
    konst_60_wire_constant <= "00000000";
    ptr_deref_55_word_offset_0 <= "0000000000000000";
    addr_of_52_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_52_final_reg_req_0;
      addr_of_52_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_52_final_reg_req_1;
      addr_of_52_final_reg_ack_1<= rack(0);
      addr_of_52_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_52_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_51_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_53,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_47_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := index_buffer(7 downto 0);
      type_cast_47_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_51_index_0_resize
    process(type_cast_47_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_47_wire;
      ov := iv(15 downto 0);
      type_cast_47_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_51_index_2_rename
    process(R_address_50_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_50_resized;
      ov(15 downto 0) := iv;
      R_address_50_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_51_index_2_resize
    process(address_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_buffer;
      ov := iv(15 downto 0);
      R_address_50_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_51_root_address_inst
    process(array_obj_ref_51_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_51_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_51_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_addr_0
    process(ptr_deref_55_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_55_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_55_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_base_resize
    process(ptr_53) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_53;
      ov := iv(15 downto 0);
      ptr_deref_55_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_gather_scatter
    process(data_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := data_buffer;
      ov(63 downto 0) := iv;
      ptr_deref_55_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_root_address_inst
    process(ptr_deref_55_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_55_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_55_root_address <= ov(15 downto 0);
      --
    end process;
    -- shared split operator group (0) : BITSEL_u8_u1_61_inst 
    ApBitsel_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= index_buffer;
      done_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= BITSEL_u8_u1_61_inst_req_0;
      BITSEL_u8_u1_61_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= BITSEL_u8_u1_61_inst_req_1;
      BITSEL_u8_u1_61_inst_ack_1 <= ackR_unguarded(0);
      ApBitsel_group_0_gI: SplitGuardInterface generic map(name => "ApBitsel_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApBitsel",
          name => "ApBitsel_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_51_index_0_scale 
    ApIntMul_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_47_resized;
      type_cast_47_scaled <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_51_index_0_scale_req_0;
      array_obj_ref_51_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_51_index_0_scale_req_1;
      array_obj_ref_51_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_1_gI: SplitGuardInterface generic map(name => "ApIntMul_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0100000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_51_index_offset 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_51_index_partial_sum_1;
      array_obj_ref_51_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_51_index_offset_req_0;
      array_obj_ref_51_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_51_index_offset_req_1;
      array_obj_ref_51_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_51_index_sum_1 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_50_scaled & type_cast_47_scaled;
      array_obj_ref_51_index_partial_sum_1 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_51_index_sum_1_req_0;
      array_obj_ref_51_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_51_index_sum_1_req_1;
      array_obj_ref_51_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared store operator group (0) : ptr_deref_55_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(15 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 8);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_55_store_0_req_0;
      ptr_deref_55_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_55_store_0_req_1;
      ptr_deref_55_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_55_word_address_0;
      data_in <= ptr_deref_55_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 16,
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(15 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end writeModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(31 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(127 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      ct_core_call_reqs : out  std_logic_vector(0 downto 0);
      ct_core_call_acks : in   std_logic_vector(0 downto 0);
      ct_core_call_data : out  std_logic_vector(175 downto 0);
      ct_core_call_tag  :  out  std_logic_vector(0 downto 0);
      ct_core_return_reqs : out  std_logic_vector(0 downto 0);
      ct_core_return_acks : in   std_logic_vector(0 downto 0);
      ct_core_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module ct_core
  component ct_core is -- 
    generic (tag_length : integer); 
    port ( -- 
      inp_d0 : in  std_logic_vector(15 downto 0);
      inp_d1 : in  std_logic_vector(15 downto 0);
      inp_d2 : in  std_logic_vector(15 downto 0);
      ker_d1 : in  std_logic_vector(15 downto 0);
      ker_d2 : in  std_logic_vector(15 downto 0);
      out_d0 : in  std_logic_vector(15 downto 0);
      out_d1 : in  std_logic_vector(15 downto 0);
      out_d2 : in  std_logic_vector(15 downto 0);
      stride : in  std_logic_vector(15 downto 0);
      padding : in  std_logic_vector(15 downto 0);
      index1 : in  std_logic_vector(7 downto 0);
      index3 : in  std_logic_vector(7 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(39 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(0 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(103 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_data : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ct_core
  signal ct_core_inp_d0 :  std_logic_vector(15 downto 0);
  signal ct_core_inp_d1 :  std_logic_vector(15 downto 0);
  signal ct_core_inp_d2 :  std_logic_vector(15 downto 0);
  signal ct_core_ker_d1 :  std_logic_vector(15 downto 0);
  signal ct_core_ker_d2 :  std_logic_vector(15 downto 0);
  signal ct_core_out_d0 :  std_logic_vector(15 downto 0);
  signal ct_core_out_d1 :  std_logic_vector(15 downto 0);
  signal ct_core_out_d2 :  std_logic_vector(15 downto 0);
  signal ct_core_stride :  std_logic_vector(15 downto 0);
  signal ct_core_padding :  std_logic_vector(15 downto 0);
  signal ct_core_index1 :  std_logic_vector(7 downto 0);
  signal ct_core_index3 :  std_logic_vector(7 downto 0);
  signal ct_core_in_args    : std_logic_vector(175 downto 0);
  signal ct_core_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ct_core_tag_out   : std_logic_vector(1 downto 0);
  signal ct_core_start_req : std_logic;
  signal ct_core_start_ack : std_logic;
  signal ct_core_fin_req   : std_logic;
  signal ct_core_fin_ack : std_logic;
  -- caller side aggregated signals for module ct_core
  signal ct_core_call_reqs: std_logic_vector(0 downto 0);
  signal ct_core_call_acks: std_logic_vector(0 downto 0);
  signal ct_core_return_reqs: std_logic_vector(0 downto 0);
  signal ct_core_return_acks: std_logic_vector(0 downto 0);
  signal ct_core_call_data: std_logic_vector(175 downto 0);
  signal ct_core_call_tag: std_logic_vector(0 downto 0);
  signal ct_core_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module readModule1
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readModule1
  signal readModule1_index :  std_logic_vector(7 downto 0);
  signal readModule1_address :  std_logic_vector(31 downto 0);
  signal readModule1_data :  std_logic_vector(63 downto 0);
  signal readModule1_in_args    : std_logic_vector(39 downto 0);
  signal readModule1_out_args   : std_logic_vector(63 downto 0);
  signal readModule1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal readModule1_tag_out   : std_logic_vector(1 downto 0);
  signal readModule1_start_req : std_logic;
  signal readModule1_start_ack : std_logic;
  signal readModule1_fin_req   : std_logic;
  signal readModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module readModule1
  signal readModule1_call_reqs: std_logic_vector(0 downto 0);
  signal readModule1_call_acks: std_logic_vector(0 downto 0);
  signal readModule1_return_reqs: std_logic_vector(0 downto 0);
  signal readModule1_return_acks: std_logic_vector(0 downto 0);
  signal readModule1_call_data: std_logic_vector(39 downto 0);
  signal readModule1_call_tag: std_logic_vector(0 downto 0);
  signal readModule1_return_data: std_logic_vector(63 downto 0);
  signal readModule1_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- declarations related to module writeModule1
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeModule1
  signal writeModule1_index :  std_logic_vector(7 downto 0);
  signal writeModule1_address :  std_logic_vector(31 downto 0);
  signal writeModule1_data :  std_logic_vector(63 downto 0);
  signal writeModule1_done :  std_logic_vector(0 downto 0);
  signal writeModule1_in_args    : std_logic_vector(103 downto 0);
  signal writeModule1_out_args   : std_logic_vector(0 downto 0);
  signal writeModule1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeModule1_tag_out   : std_logic_vector(1 downto 0);
  signal writeModule1_start_req : std_logic;
  signal writeModule1_start_ack : std_logic;
  signal writeModule1_fin_req   : std_logic;
  signal writeModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module writeModule1
  signal writeModule1_call_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_call_acks: std_logic_vector(0 downto 0);
  signal writeModule1_return_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_return_acks: std_logic_vector(0 downto 0);
  signal writeModule1_call_data: std_logic_vector(103 downto 0);
  signal writeModule1_call_tag: std_logic_vector(0 downto 0);
  signal writeModule1_return_data: std_logic_vector(0 downto 0);
  signal writeModule1_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(15 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(15 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      ct_core_call_reqs => ct_core_call_reqs(0 downto 0),
      ct_core_call_acks => ct_core_call_acks(0 downto 0),
      ct_core_call_data => ct_core_call_data(175 downto 0),
      ct_core_call_tag => ct_core_call_tag(0 downto 0),
      ct_core_return_reqs => ct_core_return_reqs(0 downto 0),
      ct_core_return_acks => ct_core_return_acks(0 downto 0),
      ct_core_return_tag => ct_core_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module ct_core
  ct_core_inp_d0 <= ct_core_in_args(175 downto 160);
  ct_core_inp_d1 <= ct_core_in_args(159 downto 144);
  ct_core_inp_d2 <= ct_core_in_args(143 downto 128);
  ct_core_ker_d1 <= ct_core_in_args(127 downto 112);
  ct_core_ker_d2 <= ct_core_in_args(111 downto 96);
  ct_core_out_d0 <= ct_core_in_args(95 downto 80);
  ct_core_out_d1 <= ct_core_in_args(79 downto 64);
  ct_core_out_d2 <= ct_core_in_args(63 downto 48);
  ct_core_stride <= ct_core_in_args(47 downto 32);
  ct_core_padding <= ct_core_in_args(31 downto 16);
  ct_core_index1 <= ct_core_in_args(15 downto 8);
  ct_core_index3 <= ct_core_in_args(7 downto 0);
  -- call arbiter for module ct_core
  ct_core_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 176,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => ct_core_call_reqs,
      call_acks => ct_core_call_acks,
      return_reqs => ct_core_return_reqs,
      return_acks => ct_core_return_acks,
      call_data  => ct_core_call_data,
      call_tag  => ct_core_call_tag,
      return_tag  => ct_core_return_tag,
      call_mtag => ct_core_tag_in,
      return_mtag => ct_core_tag_out,
      call_mreq => ct_core_start_req,
      call_mack => ct_core_start_ack,
      return_mreq => ct_core_fin_req,
      return_mack => ct_core_fin_ack,
      call_mdata => ct_core_in_args,
      clk => clk, 
      reset => reset --
    ); --
  ct_core_instance:ct_core-- 
    generic map(tag_length => 2)
    port map(-- 
      inp_d0 => ct_core_inp_d0,
      inp_d1 => ct_core_inp_d1,
      inp_d2 => ct_core_inp_d2,
      ker_d1 => ct_core_ker_d1,
      ker_d2 => ct_core_ker_d2,
      out_d0 => ct_core_out_d0,
      out_d1 => ct_core_out_d1,
      out_d2 => ct_core_out_d2,
      stride => ct_core_stride,
      padding => ct_core_padding,
      index1 => ct_core_index1,
      index3 => ct_core_index3,
      start_req => ct_core_start_req,
      start_ack => ct_core_start_ack,
      fin_req => ct_core_fin_req,
      fin_ack => ct_core_fin_ack,
      clk => clk,
      reset => reset,
      readModule1_call_reqs => readModule1_call_reqs(0 downto 0),
      readModule1_call_acks => readModule1_call_acks(0 downto 0),
      readModule1_call_data => readModule1_call_data(39 downto 0),
      readModule1_call_tag => readModule1_call_tag(0 downto 0),
      readModule1_return_reqs => readModule1_return_reqs(0 downto 0),
      readModule1_return_acks => readModule1_return_acks(0 downto 0),
      readModule1_return_data => readModule1_return_data(63 downto 0),
      readModule1_return_tag => readModule1_return_tag(0 downto 0),
      writeModule1_call_reqs => writeModule1_call_reqs(0 downto 0),
      writeModule1_call_acks => writeModule1_call_acks(0 downto 0),
      writeModule1_call_data => writeModule1_call_data(103 downto 0),
      writeModule1_call_tag => writeModule1_call_tag(0 downto 0),
      writeModule1_return_reqs => writeModule1_return_reqs(0 downto 0),
      writeModule1_return_acks => writeModule1_return_acks(0 downto 0),
      writeModule1_return_data => writeModule1_return_data(0 downto 0),
      writeModule1_return_tag => writeModule1_return_tag(0 downto 0),
      tag_in => ct_core_tag_in,
      tag_out => ct_core_tag_out-- 
    ); -- 
  -- module readModule1
  readModule1_index <= readModule1_in_args(39 downto 32);
  readModule1_address <= readModule1_in_args(31 downto 0);
  readModule1_out_args <= readModule1_data ;
  -- call arbiter for module readModule1
  readModule1_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 40,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => readModule1_call_reqs,
      call_acks => readModule1_call_acks,
      return_reqs => readModule1_return_reqs,
      return_acks => readModule1_return_acks,
      call_data  => readModule1_call_data,
      call_tag  => readModule1_call_tag,
      return_tag  => readModule1_return_tag,
      call_mtag => readModule1_tag_in,
      return_mtag => readModule1_tag_out,
      return_data =>readModule1_return_data,
      call_mreq => readModule1_start_req,
      call_mack => readModule1_start_ack,
      return_mreq => readModule1_fin_req,
      return_mack => readModule1_fin_ack,
      call_mdata => readModule1_in_args,
      return_mdata => readModule1_out_args,
      clk => clk, 
      reset => reset --
    ); --
  readModule1_instance:readModule1-- 
    generic map(tag_length => 2)
    port map(-- 
      index => readModule1_index,
      address => readModule1_address,
      data => readModule1_data,
      start_req => readModule1_start_req,
      start_ack => readModule1_start_ack,
      fin_req => readModule1_fin_req,
      fin_ack => readModule1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(31 downto 16),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      tag_in => readModule1_tag_in,
      tag_out => readModule1_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  -- module writeModule1
  writeModule1_index <= writeModule1_in_args(103 downto 96);
  writeModule1_address <= writeModule1_in_args(95 downto 64);
  writeModule1_data <= writeModule1_in_args(63 downto 0);
  writeModule1_out_args <= writeModule1_done ;
  -- call arbiter for module writeModule1
  writeModule1_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 104,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeModule1_call_reqs,
      call_acks => writeModule1_call_acks,
      return_reqs => writeModule1_return_reqs,
      return_acks => writeModule1_return_acks,
      call_data  => writeModule1_call_data,
      call_tag  => writeModule1_call_tag,
      return_tag  => writeModule1_return_tag,
      call_mtag => writeModule1_tag_in,
      return_mtag => writeModule1_tag_out,
      return_data =>writeModule1_return_data,
      call_mreq => writeModule1_start_req,
      call_mack => writeModule1_start_ack,
      return_mreq => writeModule1_fin_req,
      return_mack => writeModule1_fin_ack,
      call_mdata => writeModule1_in_args,
      return_mdata => writeModule1_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeModule1_instance:writeModule1-- 
    generic map(tag_length => 2)
    port map(-- 
      index => writeModule1_index,
      address => writeModule1_address,
      data => writeModule1_data,
      done => writeModule1_done,
      start_req => writeModule1_start_req,
      start_ack => writeModule1_start_ack,
      fin_req => writeModule1_fin_req,
      fin_ack => writeModule1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(31 downto 16),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      tag_in => writeModule1_tag_in,
      tag_out => writeModule1_tag_out-- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 2,
      addr_width => 16,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 16,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
