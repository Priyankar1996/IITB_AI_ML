-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_44_branch_req_0 : boolean;
  signal phi_stmt_46_ack_0 : boolean;
  signal phi_stmt_46_req_0 : boolean;
  signal phi_stmt_46_req_1 : boolean;
  signal n_address_280_48_buf_req_0 : boolean;
  signal n_address_280_48_buf_ack_0 : boolean;
  signal n_address_280_48_buf_req_1 : boolean;
  signal n_address_280_48_buf_ack_1 : boolean;
  signal phi_stmt_51_req_0 : boolean;
  signal phi_stmt_51_req_1 : boolean;
  signal phi_stmt_51_ack_0 : boolean;
  signal n_word_start_269_53_buf_req_0 : boolean;
  signal n_word_start_269_53_buf_ack_0 : boolean;
  signal n_word_start_269_53_buf_req_1 : boolean;
  signal n_word_start_269_53_buf_ack_1 : boolean;
  signal n_winr_209_68_buf_req_1 : boolean;
  signal n_winr_209_68_buf_ack_1 : boolean;
  signal phi_stmt_57_req_1 : boolean;
  signal phi_stmt_57_req_0 : boolean;
  signal phi_stmt_57_ack_0 : boolean;
  signal nl_start_35_59_buf_req_0 : boolean;
  signal nl_start_35_59_buf_ack_0 : boolean;
  signal nl_start_35_59_buf_req_1 : boolean;
  signal nl_start_35_59_buf_ack_1 : boolean;
  signal n_left_288_60_buf_req_0 : boolean;
  signal n_left_288_60_buf_ack_0 : boolean;
  signal n_left_288_60_buf_req_1 : boolean;
  signal n_left_288_60_buf_ack_1 : boolean;
  signal phi_stmt_61_req_1 : boolean;
  signal phi_stmt_61_req_0 : boolean;
  signal phi_stmt_61_ack_0 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal n_blk_308_65_buf_req_0 : boolean;
  signal n_blk_308_65_buf_ack_0 : boolean;
  signal n_blk_308_65_buf_req_1 : boolean;
  signal n_blk_308_65_buf_ack_1 : boolean;
  signal phi_stmt_66_req_0 : boolean;
  signal phi_stmt_66_req_1 : boolean;
  signal phi_stmt_66_ack_0 : boolean;
  signal n_winr_209_68_buf_req_0 : boolean;
  signal n_winr_209_68_buf_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_1 : boolean;
  signal phi_stmt_71_req_1 : boolean;
  signal phi_stmt_71_req_0 : boolean;
  signal phi_stmt_71_ack_0 : boolean;
  signal n_col_222_75_buf_req_0 : boolean;
  signal n_col_222_75_buf_ack_0 : boolean;
  signal n_col_222_75_buf_req_1 : boolean;
  signal n_col_222_75_buf_ack_1 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  signal n_row_234_80_buf_req_0 : boolean;
  signal n_row_234_80_buf_ack_0 : boolean;
  signal n_row_234_80_buf_req_1 : boolean;
  signal n_row_234_80_buf_ack_1 : boolean;
  signal array_obj_ref_133_index_offset_req_0 : boolean;
  signal array_obj_ref_133_index_offset_ack_0 : boolean;
  signal array_obj_ref_133_index_offset_req_1 : boolean;
  signal array_obj_ref_133_index_offset_ack_1 : boolean;
  signal addr_of_134_final_reg_req_0 : boolean;
  signal addr_of_134_final_reg_ack_0 : boolean;
  signal addr_of_134_final_reg_req_1 : boolean;
  signal addr_of_134_final_reg_ack_1 : boolean;
  signal ptr_deref_138_load_0_req_0 : boolean;
  signal ptr_deref_138_load_0_ack_0 : boolean;
  signal ptr_deref_138_load_0_req_1 : boolean;
  signal ptr_deref_138_load_0_ack_1 : boolean;
  signal slice_142_inst_req_0 : boolean;
  signal slice_142_inst_ack_0 : boolean;
  signal slice_142_inst_req_1 : boolean;
  signal slice_142_inst_ack_1 : boolean;
  signal slice_146_inst_req_0 : boolean;
  signal slice_146_inst_ack_0 : boolean;
  signal slice_146_inst_req_1 : boolean;
  signal slice_146_inst_ack_1 : boolean;
  signal slice_150_inst_req_0 : boolean;
  signal slice_150_inst_ack_0 : boolean;
  signal slice_150_inst_req_1 : boolean;
  signal slice_150_inst_ack_1 : boolean;
  signal slice_154_inst_req_0 : boolean;
  signal slice_154_inst_ack_0 : boolean;
  signal slice_154_inst_req_1 : boolean;
  signal slice_154_inst_ack_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_1 : boolean;
  signal do_while_stmt_44_branch_ack_0 : boolean;
  signal do_while_stmt_44_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__exit__
      -- CP-element group 0: 	 branch_block_stmt_26/do_while_stmt_44__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_26/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/branch_block_stmt_26__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_26/$exit
      -- CP-element group 1: 	 branch_block_stmt_26/branch_block_stmt_26__exit__
      -- CP-element group 1: 	 branch_block_stmt_26/do_while_stmt_44__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/$entry
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_26/do_while_stmt_44/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/condition_done
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_26/do_while_stmt_44/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	97 
    -- CP-element group 7: 	116 
    -- CP-element group 7: 	135 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	78 
    -- CP-element group 8: 	99 
    -- CP-element group 8: 	118 
    -- CP-element group 8: 	137 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	91 
    -- CP-element group 9: 	92 
    -- CP-element group 9: 	110 
    -- CP-element group 9: 	111 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	130 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	203 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_44_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(14) & access_T_CP_0_elements(203);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	110 
    -- CP-element group 11: 	129 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	112 
    -- CP-element group 11: 	131 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(15) & access_T_CP_0_elements(32) & access_T_CP_0_elements(51) & access_T_CP_0_elements(70) & access_T_CP_0_elements(91) & access_T_CP_0_elements(110) & access_T_CP_0_elements(129) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	94 
    -- CP-element group 12: 	113 
    -- CP-element group 12: 	132 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12: 	91 
    -- CP-element group 12: 	110 
    -- CP-element group 12: 	129 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(17) & access_T_CP_0_elements(35) & access_T_CP_0_elements(54) & access_T_CP_0_elements(73) & access_T_CP_0_elements(94) & access_T_CP_0_elements(113) & access_T_CP_0_elements(132);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: 	92 
    -- CP-element group 13: 	111 
    -- CP-element group 13: 	130 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	95 
    -- CP-element group 13: 	114 
    -- CP-element group 13: 	133 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(16) & access_T_CP_0_elements(33) & access_T_CP_0_elements(52) & access_T_CP_0_elements(71) & access_T_CP_0_elements(92) & access_T_CP_0_elements(111) & access_T_CP_0_elements(130);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	96 
    -- CP-element group 14: 	115 
    -- CP-element group 14: 	134 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(56) & access_T_CP_0_elements(75) & access_T_CP_0_elements(96) & access_T_CP_0_elements(115) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	151 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (15) 
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/req
      -- 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(18), ack => array_obj_ref_133_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_trigger
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req_ps
      -- 
    phi_stmt_46_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => phi_stmt_46_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req_ps
      -- 
    phi_stmt_46_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_46_req_1); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack_ps
      -- 
    phi_stmt_46_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_46_ack_0, ack => access_T_CP_0_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Sample/req
      -- 
    req_63_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_63_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => n_address_280_48_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_update_start_
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Update/req
      -- 
    req_68_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_68_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(25), ack => n_address_280_48_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Sample/ack
      -- 
    ack_64_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_48_buf_ack_0, ack => access_T_CP_0_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_48_Update/ack
      -- 
    ack_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_48_buf_ack_1, ack => access_T_CP_0_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_update_start_
      -- 
    -- Element group access_T_CP_0_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_update_completed__ps
      -- 
    access_T_CP_0_elements(30) <= access_T_CP_0_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_50_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(29), ack => access_T_CP_0_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start_
      -- 
    access_T_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	191 
    -- CP-element group 33: 	177 
    -- CP-element group 33: 	184 
    -- CP-element group 33: 	198 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start_
      -- 
    access_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(191) & access_T_CP_0_elements(177) & access_T_CP_0_elements(184) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start__ps
      -- 
    access_T_CP_0_elements(34) <= access_T_CP_0_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	196 
    -- CP-element group 37: 	175 
    -- CP-element group 37: 	182 
    -- CP-element group 37: 	189 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_trigger
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req_ps
      -- 
    phi_stmt_51_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(39), ack => phi_stmt_51_req_0); -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req_ps
      -- 
    phi_stmt_51_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_51_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack_ps
      -- 
    phi_stmt_51_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_51_ack_0, ack => access_T_CP_0_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Sample/req
      -- 
    req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => n_word_start_269_53_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_update_start_
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Update/req
      -- 
    req_112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(44), ack => n_word_start_269_53_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Sample/ack
      -- 
    ack_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_53_buf_ack_0, ack => access_T_CP_0_elements(45)); -- 
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_53_Update/ack
      -- 
    ack_113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_53_buf_ack_1, ack => access_T_CP_0_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_update_start_
      -- 
    -- Element group access_T_CP_0_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_update_completed__ps
      -- 
    access_T_CP_0_elements(49) <= access_T_CP_0_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_56_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(48), ack => access_T_CP_0_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start_
      -- 
    access_T_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	56 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start_
      -- 
    access_T_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(56);
      gj_access_T_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start__ps
      -- 
    access_T_CP_0_elements(53) <= access_T_CP_0_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start__ps
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_trigger
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req_ps
      -- 
    phi_stmt_57_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(58), ack => phi_stmt_57_req_1); -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_trigger
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req_ps
      -- 
    phi_stmt_57_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => phi_stmt_57_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack_ps
      -- 
    phi_stmt_57_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_57_ack_0, ack => access_T_CP_0_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/req
      -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => nl_start_35_59_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start_
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/req
      -- 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(63), ack => nl_start_35_59_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_0, ack => access_T_CP_0_elements(64)); -- 
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_1, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(66), ack => n_left_288_60_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start_
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(67), ack => n_left_288_60_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_0, ack => access_T_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_1, ack => access_T_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start_
      -- 
    access_T_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	191 
    -- CP-element group 71: 	184 
    -- CP-element group 71: 	198 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start_
      -- 
    access_T_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(191) & access_T_CP_0_elements(184) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start__ps
      -- 
    access_T_CP_0_elements(72) <= access_T_CP_0_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start__ps
      -- 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	196 
    -- CP-element group 75: 	182 
    -- CP-element group 75: 	189 
    -- CP-element group 75: 	14 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_trigger
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req_ps
      -- 
    phi_stmt_61_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(77), ack => phi_stmt_61_req_1); -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req_ps
      -- 
    phi_stmt_61_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_61_req_0); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack_ps
      -- 
    phi_stmt_61_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_61_ack_0, ack => access_T_CP_0_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/rr
      -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => type_cast_64_inst_req_0); -- 
    access_T_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(85);
      gj_access_T_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start_
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/cr
      -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(84), ack => type_cast_64_inst_req_1); -- 
    access_T_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(82) & access_T_CP_0_elements(86);
      gj_access_T_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => access_T_CP_0_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/req
      -- 
    req_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(87), ack => n_blk_308_65_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start_
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/req
      -- 
    req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => n_blk_308_65_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/ack
      -- 
    ack_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_0, ack => access_T_CP_0_elements(89)); -- 
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/ack
      -- 
    ack_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_1, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	9 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	12 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	11 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start_
      -- 
    access_T_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	9 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	96 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	13 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start_
      -- 
    access_T_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(96);
      gj_access_T_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	11 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start__ps
      -- 
    access_T_CP_0_elements(93) <= access_T_CP_0_elements(11);
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	12 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	13 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start__ps
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(13);
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	14 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	92 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	7 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_trigger
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(7);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req_ps
      -- 
    phi_stmt_66_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => phi_stmt_66_req_0); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	8 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(8);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req_ps
      -- 
    phi_stmt_66_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_66_req_1); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack_ps
      -- 
    phi_stmt_66_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_66_ack_0, ack => access_T_CP_0_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_start__ps
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/req
      -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(102), ack => n_winr_209_68_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/req
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_start__ps
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_start_
      -- 
    req_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(103), ack => n_winr_209_68_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_68_buf_ack_0, ack => access_T_CP_0_elements(104)); -- 
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/ack
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_completed__ps
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_completed_
      -- 
    ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_68_buf_ack_1, ack => access_T_CP_0_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_start_
      -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_completed__ps
      -- 
    access_T_CP_0_elements(108) <= access_T_CP_0_elements(109);
    -- CP-element group 109:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	108 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(107), ack => access_T_CP_0_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	9 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	12 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	11 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start_
      -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	115 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	13 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start_
      -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(115);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	11 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start__ps
      -- 
    access_T_CP_0_elements(112) <= access_T_CP_0_elements(11);
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	12 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	13 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(13);
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	14 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	111 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	7 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_trigger
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(7);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req_ps
      -- 
    phi_stmt_71_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_71_req_1); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	8 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_trigger
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(8);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req_ps
      -- 
    phi_stmt_71_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_71_req_0); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack_ps
      -- 
    phi_stmt_71_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_71_ack_0, ack => access_T_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_start_
      -- 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_completed__ps
      -- 
    access_T_CP_0_elements(123) <= access_T_CP_0_elements(124);
    -- CP-element group 124:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(124) is a control-delay.
    cp_element_124_delay: control_delay_element  generic map(name => " 124_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(122), ack => access_T_CP_0_elements(124), clk => clk, reset =>reset);
    -- CP-element group 125:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/req
      -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => n_col_222_75_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_start_
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/req
      -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(126), ack => n_col_222_75_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/ack
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_75_buf_ack_0, ack => access_T_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_75_buf_ack_1, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	12 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	11 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start_
      -- 
    access_T_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	9 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	134 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	13 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start_
      -- 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	11 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start__ps
      -- 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(11);
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	12 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start__ps
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(13);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	130 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req_ps
      -- 
    phi_stmt_76_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_76_req_1); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_trigger
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req_ps
      -- 
    phi_stmt_76_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_76_req_0); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack_ps
      -- 
    phi_stmt_76_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_start_
      -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_completed__ps
      -- 
    access_T_CP_0_elements(142) <= access_T_CP_0_elements(143);
    -- CP-element group 143:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(141), ack => access_T_CP_0_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/req
      -- 
    req_355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(144), ack => n_row_234_80_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (4) 
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_start_
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/req
      -- 
    req_360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(145), ack => n_row_234_80_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/ack
      -- 
    ack_356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_80_buf_ack_0, ack => access_T_CP_0_elements(146)); -- 
    -- CP-element group 147:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_completed__ps
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/ack
      -- 
    ack_361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_80_buf_ack_1, ack => access_T_CP_0_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_134_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_start_
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_134_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/req
      -- 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_133_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	18 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/ack
      -- 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_ack
      -- 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: 	148 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/rr
      -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_138_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	173 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	169 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_start_
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/cr
      -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_138_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(173) & access_T_CP_0_elements(161) & access_T_CP_0_elements(165) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: 	149 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158: 	167 
    -- CP-element group 158: 	171 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_ack
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/rr
      -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_142_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_start_
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/cr
      -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_142_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/rr
      -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_146_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_start_
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/cr
      -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_146_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	156 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/rr
      -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_150_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_start_
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/cr
      -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_150_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	156 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/rr
      -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_154_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_start_
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/cr
      -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_154_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: 	156 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	37 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_156_delayed_14_0_156_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_start_
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/req
      -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_156_delayed_14_0_156_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	33 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	162 
    -- CP-element group 179: 	178 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_160_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(162) & access_T_CP_0_elements(178) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	160 
    -- CP-element group 180: 	176 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_start_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_160_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	37 
    -- CP-element group 182: 	75 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_160_delayed_14_0_163_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_start_
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_160_delayed_14_0_163_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	33 
    -- CP-element group 184: 	71 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	166 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	181 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_167_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(166) & access_T_CP_0_elements(185) & access_T_CP_0_elements(181) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: 	164 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/req
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_start_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$exit
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_167_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_completed_
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	37 
    -- CP-element group 189: 	75 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_164_delayed_14_0_170_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_start_
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/req
      -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_164_delayed_14_0_170_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	33 
    -- CP-element group 191: 	71 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	170 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/req
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_174_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(192) & access_T_CP_0_elements(188) & access_T_CP_0_elements(170) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	168 
    -- CP-element group 194: 	190 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_start_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/req
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_174_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	37 
    -- CP-element group 196: 	75 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/req
      -- 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_168_delayed_14_0_177_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_start_
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/req
      -- 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_168_delayed_14_0_177_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	33 
    -- CP-element group 198: 	71 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/ack
      -- 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	174 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_181_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(195) & access_T_CP_0_elements(174) & access_T_CP_0_elements(199) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	197 
    -- CP-element group 201: 	172 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_start_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/req
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_181_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	179 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	151 
    -- CP-element group 204: 	12 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$exit
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(151) & access_T_CP_0_elements(12) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/ack
      -- 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_26/do_while_stmt_44/$exit
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_44_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_44_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_46_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(19);
      access_T_CP_0_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(27);
      access_T_CP_0_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(30);
      access_T_CP_0_elements(22) <= phi_mux_reqs(1);
      phi_stmt_46_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_46_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(17), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(18), 
          phi_mux_ack => access_T_CP_0_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_51_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(38);
      access_T_CP_0_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(46);
      access_T_CP_0_elements(39) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(49);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_51_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_51_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(34), 
          phi_sample_ack => access_T_CP_0_elements(35), 
          phi_update_req => access_T_CP_0_elements(36), 
          phi_update_ack => access_T_CP_0_elements(37), 
          phi_mux_ack => access_T_CP_0_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_57_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(59);
      access_T_CP_0_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(64);
      access_T_CP_0_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(65);
      access_T_CP_0_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(57);
      access_T_CP_0_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(68);
      access_T_CP_0_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(69);
      access_T_CP_0_elements(58) <= phi_mux_reqs(1);
      phi_stmt_57_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_57_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(53), 
          phi_sample_ack => access_T_CP_0_elements(54), 
          phi_update_req => access_T_CP_0_elements(55), 
          phi_update_ack => access_T_CP_0_elements(56), 
          phi_mux_ack => access_T_CP_0_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_61_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(85);
      access_T_CP_0_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(86);
      access_T_CP_0_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(76);
      access_T_CP_0_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(77) <= phi_mux_reqs(1);
      phi_stmt_61_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_61_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(72), 
          phi_sample_ack => access_T_CP_0_elements(73), 
          phi_update_req => access_T_CP_0_elements(74), 
          phi_update_ack => access_T_CP_0_elements(75), 
          phi_mux_ack => access_T_CP_0_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_66_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(97);
      access_T_CP_0_elements(102)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(103)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(105);
      access_T_CP_0_elements(98) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(106)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(106);
      access_T_CP_0_elements(107)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(108);
      access_T_CP_0_elements(100) <= phi_mux_reqs(1);
      phi_stmt_66_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_66_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(93), 
          phi_sample_ack => access_T_CP_0_elements(94), 
          phi_update_req => access_T_CP_0_elements(95), 
          phi_update_ack => access_T_CP_0_elements(96), 
          phi_mux_ack => access_T_CP_0_elements(101), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_71_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(121)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(121);
      access_T_CP_0_elements(122)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(123);
      access_T_CP_0_elements(119) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(125)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(126)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(128);
      access_T_CP_0_elements(117) <= phi_mux_reqs(1);
      phi_stmt_71_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_71_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(112), 
          phi_sample_ack => access_T_CP_0_elements(113), 
          phi_update_req => access_T_CP_0_elements(114), 
          phi_update_ack => access_T_CP_0_elements(115), 
          phi_mux_ack => access_T_CP_0_elements(120), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_76_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(140);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(138) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(147);
      access_T_CP_0_elements(136) <= phi_mux_reqs(1);
      phi_stmt_76_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_76_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(131), 
          phi_sample_ack => access_T_CP_0_elements(132), 
          phi_update_req => access_T_CP_0_elements(133), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_125_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_205_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_218_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_231_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_241_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_293_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_278_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_107_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_114_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_213_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_227_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_228_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_94_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_260_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_103_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_110_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_117_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_90_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_97_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_274_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_240_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_30_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_249_wire : std_logic_vector(31 downto 0);
    signal MUX_206_wire : std_logic_vector(15 downto 0);
    signal MUX_219_wire : std_logic_vector(15 downto 0);
    signal MUX_300_wire : std_logic_vector(15 downto 0);
    signal MUX_306_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_312_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_118_wire : std_logic_vector(0 downto 0);
    signal R_address_132_resized : std_logic_vector(13 downto 0);
    signal R_address_132_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_286_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_298_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_106_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_113_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_295_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_93_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_303_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_39_wire : std_logic_vector(0 downto 0);
    signal address_46 : std_logic_vector(63 downto 0);
    signal array_obj_ref_133_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_root_address : std_logic_vector(13 downto 0);
    signal c1_156_delayed_14_0_158 : std_logic_vector(0 downto 0);
    signal c1_86 : std_logic_vector(0 downto 0);
    signal c2_160_delayed_14_0_165 : std_logic_vector(0 downto 0);
    signal c2_99 : std_logic_vector(0 downto 0);
    signal c3_120 : std_logic_vector(0 downto 0);
    signal c3_164_delayed_14_0_172 : std_logic_vector(0 downto 0);
    signal c4_128 : std_logic_vector(0 downto 0);
    signal c4_168_delayed_14_0_179 : std_logic_vector(0 downto 0);
    signal col_71 : std_logic_vector(15 downto 0);
    signal col_done_198 : std_logic_vector(0 downto 0);
    signal fetch_addr_135 : std_logic_vector(31 downto 0);
    signal flag1_188 : std_logic_vector(0 downto 0);
    signal fn_blk_43 : std_logic_vector(15 downto 0);
    signal konst_102_wire_constant : std_logic_vector(1 downto 0);
    signal konst_105_wire_constant : std_logic_vector(15 downto 0);
    signal konst_109_wire_constant : std_logic_vector(1 downto 0);
    signal konst_112_wire_constant : std_logic_vector(15 downto 0);
    signal konst_116_wire_constant : std_logic_vector(1 downto 0);
    signal konst_126_wire_constant : std_logic_vector(15 downto 0);
    signal konst_202_wire_constant : std_logic_vector(15 downto 0);
    signal konst_204_wire_constant : std_logic_vector(15 downto 0);
    signal konst_215_wire_constant : std_logic_vector(15 downto 0);
    signal konst_217_wire_constant : std_logic_vector(15 downto 0);
    signal konst_230_wire_constant : std_logic_vector(15 downto 0);
    signal konst_259_wire_constant : std_logic_vector(31 downto 0);
    signal konst_267_wire_constant : std_logic_vector(1 downto 0);
    signal konst_273_wire_constant : std_logic_vector(31 downto 0);
    signal konst_277_wire_constant : std_logic_vector(63 downto 0);
    signal konst_294_wire_constant : std_logic_vector(15 downto 0);
    signal konst_296_wire_constant : std_logic_vector(15 downto 0);
    signal konst_302_wire_constant : std_logic_vector(15 downto 0);
    signal konst_305_wire_constant : std_logic_vector(15 downto 0);
    signal konst_38_wire_constant : std_logic_vector(15 downto 0);
    signal konst_41_wire_constant : std_logic_vector(15 downto 0);
    signal konst_84_wire_constant : std_logic_vector(1 downto 0);
    signal konst_89_wire_constant : std_logic_vector(1 downto 0);
    signal konst_92_wire_constant : std_logic_vector(15 downto 0);
    signal konst_96_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_32 : std_logic_vector(31 downto 0);
    signal n_address_280 : std_logic_vector(63 downto 0);
    signal n_address_280_48_buffered : std_logic_vector(63 downto 0);
    signal n_blk_308 : std_logic_vector(15 downto 0);
    signal n_blk_308_65_buffered : std_logic_vector(15 downto 0);
    signal n_col_222 : std_logic_vector(15 downto 0);
    signal n_col_222_75_buffered : std_logic_vector(15 downto 0);
    signal n_left_288 : std_logic_vector(15 downto 0);
    signal n_left_288_60_buffered : std_logic_vector(15 downto 0);
    signal n_row_234 : std_logic_vector(15 downto 0);
    signal n_row_234_80_buffered : std_logic_vector(15 downto 0);
    signal n_winr_209 : std_logic_vector(15 downto 0);
    signal n_winr_209_68_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_269 : std_logic_vector(1 downto 0);
    signal n_word_start_269_53_buffered : std_logic_vector(1 downto 0);
    signal na1_244 : std_logic_vector(31 downto 0);
    signal na2_251 : std_logic_vector(31 downto 0);
    signal na3_256 : std_logic_vector(31 downto 0);
    signal na4_262 : std_logic_vector(15 downto 0);
    signal nl_start_35 : std_logic_vector(15 downto 0);
    signal nl_start_35_59_buffered : std_logic_vector(15 downto 0);
    signal num_blk_61 : std_logic_vector(15 downto 0);
    signal num_left_57 : std_logic_vector(15 downto 0);
    signal ptr_deref_138_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_138_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_76 : std_logic_vector(15 downto 0);
    signal type_cast_124_wire : std_logic_vector(15 downto 0);
    signal type_cast_248_wire : std_logic_vector(31 downto 0);
    signal type_cast_266_wire : std_logic_vector(1 downto 0);
    signal type_cast_275_wire : std_logic_vector(63 downto 0);
    signal type_cast_50_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_56_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_64_wire : std_logic_vector(15 downto 0);
    signal type_cast_70_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_74_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(15 downto 0);
    signal w1_143 : std_logic_vector(15 downto 0);
    signal w2_147 : std_logic_vector(15 downto 0);
    signal w3_151 : std_logic_vector(15 downto 0);
    signal w4_155 : std_logic_vector(15 downto 0);
    signal winr_66 : std_logic_vector(15 downto 0);
    signal winr_done_193 : std_logic_vector(0 downto 0);
    signal word_read_139 : std_logic_vector(63 downto 0);
    signal word_start_51 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_133_constant_part_of_offset <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_133_resized_base_address <= "00000000000000";
    konst_102_wire_constant <= "00";
    konst_105_wire_constant <= "0000000000000010";
    konst_109_wire_constant <= "01";
    konst_112_wire_constant <= "0000000000000001";
    konst_116_wire_constant <= "10";
    konst_126_wire_constant <= "0000000000000011";
    konst_202_wire_constant <= "0000000000000000";
    konst_204_wire_constant <= "0000000000000001";
    konst_215_wire_constant <= "0000000000000000";
    konst_217_wire_constant <= "0000000000000001";
    konst_230_wire_constant <= "0000000000000001";
    konst_259_wire_constant <= "00000000000000000000000000000011";
    konst_267_wire_constant <= "00";
    konst_273_wire_constant <= "00000000000000000000000000000010";
    konst_277_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_294_wire_constant <= "0000000000000100";
    konst_296_wire_constant <= "0000000000000100";
    konst_302_wire_constant <= "0000000000000100";
    konst_305_wire_constant <= "0000000000000100";
    konst_38_wire_constant <= "0000000000000100";
    konst_41_wire_constant <= "0000000000000100";
    konst_84_wire_constant <= "00";
    konst_89_wire_constant <= "00";
    konst_92_wire_constant <= "0000000000000001";
    konst_96_wire_constant <= "01";
    ptr_deref_138_word_offset_0 <= "00000000000000";
    type_cast_50_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_56_wire_constant <= "00";
    type_cast_70_wire_constant <= "0000000000000000";
    type_cast_74_wire_constant <= "0000000000000000";
    type_cast_79_wire_constant <= "0000000000000000";
    phi_stmt_46: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address_280_48_buffered & type_cast_50_wire_constant;
      req <= phi_stmt_46_req_0 & phi_stmt_46_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_46",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_46_ack_0,
          idata => idata,
          odata => address_46,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_46
    phi_stmt_51: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_word_start_269_53_buffered & type_cast_56_wire_constant;
      req <= phi_stmt_51_req_0 & phi_stmt_51_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_51",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_51_ack_0,
          idata => idata,
          odata => word_start_51,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_51
    phi_stmt_57: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nl_start_35_59_buffered & n_left_288_60_buffered;
      req <= phi_stmt_57_req_0 & phi_stmt_57_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_57",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_57_ack_0,
          idata => idata,
          odata => num_left_57,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_57
    phi_stmt_61: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_64_wire & n_blk_308_65_buffered;
      req <= phi_stmt_61_req_0 & phi_stmt_61_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_61",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_61_ack_0,
          idata => idata,
          odata => num_blk_61,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_61
    phi_stmt_66: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_winr_209_68_buffered & type_cast_70_wire_constant;
      req <= phi_stmt_66_req_0 & phi_stmt_66_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_66",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_66_ack_0,
          idata => idata,
          odata => winr_66,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_66
    phi_stmt_71: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_74_wire_constant & n_col_222_75_buffered;
      req <= phi_stmt_71_req_0 & phi_stmt_71_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_71",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_71_ack_0,
          idata => idata,
          odata => col_71,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_71
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_79_wire_constant & n_row_234_80_buffered;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => row_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    -- flow-through select operator MUX_206_inst
    MUX_206_wire <= konst_202_wire_constant when (winr_done_193(0) /=  '0') else ADD_u16_u16_205_wire;
    -- flow-through select operator MUX_208_inst
    n_winr_209 <= MUX_206_wire when (flag1_188(0) /=  '0') else winr_66;
    -- flow-through select operator MUX_219_inst
    MUX_219_wire <= konst_215_wire_constant when (col_done_198(0) /=  '0') else ADD_u16_u16_218_wire;
    -- flow-through select operator MUX_221_inst
    n_col_222 <= MUX_219_wire when (AND_u1_u1_213_wire(0) /=  '0') else col_71;
    -- flow-through select operator MUX_233_inst
    n_row_234 <= ADD_u16_u16_231_wire when (AND_u1_u1_228_wire(0) /=  '0') else row_76;
    -- flow-through select operator MUX_268_inst
    n_word_start_269 <= type_cast_266_wire when (flag1_188(0) /=  '0') else konst_267_wire_constant;
    -- flow-through select operator MUX_279_inst
    n_address_280 <= type_cast_275_wire when (flag1_188(0) /=  '0') else ADD_u64_u64_278_wire;
    -- flow-through select operator MUX_287_inst
    n_left_288 <= nl_start_35 when (flag1_188(0) /=  '0') else SUB_u16_u16_286_wire;
    -- flow-through select operator MUX_300_inst
    MUX_300_wire <= SUB_u16_u16_298_wire when (UGT_u16_u1_295_wire(0) /=  '0') else fn_blk_43;
    -- flow-through select operator MUX_306_inst
    MUX_306_wire <= n_left_288 when (ULT_u16_u1_303_wire(0) /=  '0') else konst_305_wire_constant;
    -- flow-through select operator MUX_307_inst
    n_blk_308 <= MUX_300_wire when (flag1_188(0) /=  '0') else MUX_306_wire;
    -- flow-through select operator MUX_42_inst
    fn_blk_43 <= num_cont_buffer when (ULT_u16_u1_39_wire(0) /=  '0') else konst_41_wire_constant;
    slice_142_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_142_inst_req_0;
      slice_142_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_142_inst_req_1;
      slice_142_inst_ack_1<= update_ack(0);
      slice_142_inst: SliceSplitProtocol generic map(name => "slice_142_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w1_143, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_146_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_146_inst_req_0;
      slice_146_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_146_inst_req_1;
      slice_146_inst_ack_1<= update_ack(0);
      slice_146_inst: SliceSplitProtocol generic map(name => "slice_146_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w2_147, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_150_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_150_inst_req_0;
      slice_150_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_150_inst_req_1;
      slice_150_inst_ack_1<= update_ack(0);
      slice_150_inst: SliceSplitProtocol generic map(name => "slice_150_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w3_151, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_154_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_154_inst_req_0;
      slice_154_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_154_inst_req_1;
      slice_154_inst_ack_1<= update_ack(0);
      slice_154_inst: SliceSplitProtocol generic map(name => "slice_154_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w4_155, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_c1_156_delayed_14_0_156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_156_delayed_14_0_156_inst_req_0;
      W_c1_156_delayed_14_0_156_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_156_delayed_14_0_156_inst_req_1;
      W_c1_156_delayed_14_0_156_inst_ack_1<= rack(0);
      W_c1_156_delayed_14_0_156_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_156_delayed_14_0_156_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_156_delayed_14_0_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c2_160_delayed_14_0_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_160_delayed_14_0_163_inst_req_0;
      W_c2_160_delayed_14_0_163_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_160_delayed_14_0_163_inst_req_1;
      W_c2_160_delayed_14_0_163_inst_ack_1<= rack(0);
      W_c2_160_delayed_14_0_163_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_160_delayed_14_0_163_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_160_delayed_14_0_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c3_164_delayed_14_0_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_164_delayed_14_0_170_inst_req_0;
      W_c3_164_delayed_14_0_170_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_164_delayed_14_0_170_inst_req_1;
      W_c3_164_delayed_14_0_170_inst_ack_1<= rack(0);
      W_c3_164_delayed_14_0_170_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_164_delayed_14_0_170_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_164_delayed_14_0_172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c4_168_delayed_14_0_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_168_delayed_14_0_177_inst_req_0;
      W_c4_168_delayed_14_0_177_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_168_delayed_14_0_177_inst_req_1;
      W_c4_168_delayed_14_0_177_inst_ack_1<= rack(0);
      W_c4_168_delayed_14_0_177_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_168_delayed_14_0_177_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_168_delayed_14_0_179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nl_start_33_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_35 <= tmp_var; -- 
    end process;
    addr_of_134_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_134_final_reg_req_0;
      addr_of_134_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_134_final_reg_req_1;
      addr_of_134_final_reg_ack_1<= rack(0);
      addr_of_134_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_134_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_133_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_280_48_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_280_48_buf_req_0;
      n_address_280_48_buf_ack_0<= wack(0);
      rreq(0) <= n_address_280_48_buf_req_1;
      n_address_280_48_buf_ack_1<= rack(0);
      n_address_280_48_buf : InterlockBuffer generic map ( -- 
        name => "n_address_280_48_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_280_48_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_blk_308_65_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_308_65_buf_req_0;
      n_blk_308_65_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_308_65_buf_req_1;
      n_blk_308_65_buf_ack_1<= rack(0);
      n_blk_308_65_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_308_65_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_308_65_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_222_75_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_222_75_buf_req_0;
      n_col_222_75_buf_ack_0<= wack(0);
      rreq(0) <= n_col_222_75_buf_req_1;
      n_col_222_75_buf_ack_1<= rack(0);
      n_col_222_75_buf : InterlockBuffer generic map ( -- 
        name => "n_col_222_75_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_222_75_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_left_288_60_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_288_60_buf_req_0;
      n_left_288_60_buf_ack_0<= wack(0);
      rreq(0) <= n_left_288_60_buf_req_1;
      n_left_288_60_buf_ack_1<= rack(0);
      n_left_288_60_buf : InterlockBuffer generic map ( -- 
        name => "n_left_288_60_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_288_60_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_234_80_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_234_80_buf_req_0;
      n_row_234_80_buf_ack_0<= wack(0);
      rreq(0) <= n_row_234_80_buf_req_1;
      n_row_234_80_buf_ack_1<= rack(0);
      n_row_234_80_buf : InterlockBuffer generic map ( -- 
        name => "n_row_234_80_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_234_80_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_winr_209_68_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_209_68_buf_req_0;
      n_winr_209_68_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_209_68_buf_req_1;
      n_winr_209_68_buf_ack_1<= rack(0);
      n_winr_209_68_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_209_68_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_209_68_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_word_start_269_53_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_269_53_buf_req_0;
      n_word_start_269_53_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_269_53_buf_req_1;
      n_word_start_269_53_buf_ack_1<= rack(0);
      n_word_start_269_53_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_269_53_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_269_53_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nl_start_35_59_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_35_59_buf_req_0;
      nl_start_35_59_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_35_59_buf_req_1;
      nl_start_35_59_buf_ack_1<= rack(0);
      nl_start_35_59_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_35_59_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_35_59_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_124_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_51(1 downto 0);
      type_cast_124_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_243_inst
    process(MUL_u16_u16_242_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_242_wire(15 downto 0);
      na1_244 <= tmp_var; -- 
    end process;
    -- interlock type_cast_248_inst
    process(n_winr_209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_209(15 downto 0);
      type_cast_248_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_250_inst
    process(MUL_u32_u32_249_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_249_wire(31 downto 0);
      na2_251 <= tmp_var; -- 
    end process;
    -- interlock type_cast_261_inst
    process(AND_u32_u32_260_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_260_wire(15 downto 0);
      na4_262 <= tmp_var; -- 
    end process;
    -- interlock type_cast_266_inst
    process(na4_262) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_262(1 downto 0);
      type_cast_266_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_275_inst
    process(LSHR_u32_u32_274_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_274_wire(31 downto 0);
      type_cast_275_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_31_inst
    process(MUL_u16_u16_30_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_30_wire(15 downto 0);
      m_factor_32 <= tmp_var; -- 
    end process;
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_43,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_64_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_133_index_1_rename
    process(R_address_132_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_132_resized;
      ov(13 downto 0) := iv;
      R_address_132_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_index_1_resize
    process(address_46) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_46;
      ov := iv(13 downto 0);
      R_address_132_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_root_address_inst
    process(array_obj_ref_133_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_133_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_133_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_addr_0
    process(ptr_deref_138_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_base_resize
    process(fetch_addr_135) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_135;
      ov := iv(13 downto 0);
      ptr_deref_138_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_gather_scatter
    process(ptr_deref_138_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_data_0;
      ov(63 downto 0) := iv;
      word_read_139 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_root_address_inst
    process(ptr_deref_138_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_44_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_312_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_44_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_44_branch_req_0,
          ack0 => do_while_stmt_44_branch_ack_0,
          ack1 => do_while_stmt_44_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_125_inst
    process(num_blk_61, type_cast_124_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_61, type_cast_124_wire, tmp_var);
      ADD_u16_u16_125_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_205_inst
    process(winr_66) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_66, konst_204_wire_constant, tmp_var);
      ADD_u16_u16_205_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_218_inst
    process(col_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_71, konst_217_wire_constant, tmp_var);
      ADD_u16_u16_218_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_231_inst
    process(row_76) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_76, konst_230_wire_constant, tmp_var);
      ADD_u16_u16_231_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_241_inst
    process(n_col_222, MUL_u16_u16_240_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_222, MUL_u16_u16_240_wire, tmp_var);
      ADD_u16_u16_241_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_293_inst
    process(fn_blk_43, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_43, na4_262, tmp_var);
      ADD_u16_u16_293_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_255_inst
    process(na1_244, na2_251) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_244, na2_251, tmp_var);
      na3_256 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_278_inst
    process(address_46) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_46, konst_277_wire_constant, tmp_var);
      ADD_u64_u64_278_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_107_inst
    process(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire, tmp_var);
      AND_u1_u1_107_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_114_inst
    process(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire, tmp_var);
      AND_u1_u1_114_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_213_inst
    process(winr_done_193, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, flag1_188, tmp_var);
      AND_u1_u1_213_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_227_inst
    process(col_done_198, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_198, flag1_188, tmp_var);
      AND_u1_u1_227_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_228_inst
    process(winr_done_193, AND_u1_u1_227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, AND_u1_u1_227_wire, tmp_var);
      AND_u1_u1_228_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_94_inst
    process(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire, tmp_var);
      AND_u1_u1_94_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_260_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_256, konst_259_wire_constant, tmp_var);
      AND_u32_u32_260_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_187_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_57, num_blk_61, tmp_var);
      flag1_188 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_192_inst
    process(winr_66, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_66, rk1_buffer, tmp_var);
      winr_done_193 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_197_inst
    process(col_71, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_71, col1_buffer, tmp_var);
      col_done_198 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_103_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_102_wire_constant, tmp_var);
      EQ_u2_u1_103_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_110_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_109_wire_constant, tmp_var);
      EQ_u2_u1_110_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_117_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_116_wire_constant, tmp_var);
      EQ_u2_u1_117_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_85_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_84_wire_constant, tmp_var);
      c1_86 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_90_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_89_wire_constant, tmp_var);
      EQ_u2_u1_90_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_97_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_96_wire_constant, tmp_var);
      EQ_u2_u1_97_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_274_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_256, konst_273_wire_constant, tmp_var);
      LSHR_u32_u32_274_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_240_inst
    process(ct_buffer, n_row_234) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_234, tmp_var);
      MUL_u16_u16_240_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_242_inst
    process(chl_in_buffer, ADD_u16_u16_241_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_241_wire, tmp_var);
      MUL_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_30_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_30_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_249_inst
    process(m_factor_32, type_cast_248_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_32, type_cast_248_wire, tmp_var);
      MUL_u32_u32_249_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u16_u1_312_inst
    process(n_row_234, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_234, row1_buffer, tmp_var);
      NEQ_u16_u1_312_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_118_inst
    process(AND_u1_u1_114_wire, EQ_u2_u1_117_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_114_wire, EQ_u2_u1_117_wire, tmp_var);
      OR_u1_u1_118_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_119_inst
    process(AND_u1_u1_107_wire, OR_u1_u1_118_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_107_wire, OR_u1_u1_118_wire, tmp_var);
      c3_120 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_98_inst
    process(AND_u1_u1_94_wire, EQ_u2_u1_97_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_94_wire, EQ_u2_u1_97_wire, tmp_var);
      c2_99 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_286_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_57, num_blk_61, tmp_var);
      SUB_u16_u16_286_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_298_inst
    process(konst_296_wire_constant, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_296_wire_constant, na4_262, tmp_var);
      SUB_u16_u16_298_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_106_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_105_wire_constant, tmp_var);
      UGT_u16_u1_106_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_113_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_112_wire_constant, tmp_var);
      UGT_u16_u1_113_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_127_inst
    process(ADD_u16_u16_125_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_125_wire, konst_126_wire_constant, tmp_var);
      c4_128 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_295_inst
    process(ADD_u16_u16_293_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_293_wire, konst_294_wire_constant, tmp_var);
      UGT_u16_u1_295_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_93_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_92_wire_constant, tmp_var);
      UGT_u16_u1_93_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_303_inst
    process(n_left_288) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_288, konst_302_wire_constant, tmp_var);
      ULT_u16_u1_303_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_39_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_38_wire_constant, tmp_var);
      ULT_u16_u1_39_wire <= tmp_var; --
    end process;
    -- shared split operator group (42) : array_obj_ref_133_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_132_scaled;
      array_obj_ref_133_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_133_index_offset_req_0;
      array_obj_ref_133_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_133_index_offset_req_1;
      array_obj_ref_133_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared load operator group (0) : ptr_deref_138_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_138_load_0_req_0;
      ptr_deref_138_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_138_load_0_req_1;
      ptr_deref_138_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_138_word_address_0;
      ptr_deref_138_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_174_inst WPIPE_input_pipe1_167_inst WPIPE_input_pipe1_160_inst WPIPE_input_pipe1_181_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_174_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_167_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_160_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_0;
      WPIPE_input_pipe1_174_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_167_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_160_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_174_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_167_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_160_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_1;
      WPIPE_input_pipe1_174_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_167_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_160_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c4_168_delayed_14_0_179(0);
      guard_vector(1)  <= c1_156_delayed_14_0_158(0);
      guard_vector(2)  <= c2_160_delayed_14_0_165(0);
      guard_vector(3)  <= c3_164_delayed_14_0_172(0);
      data_in <= w3_151 & w2_147 & w1_143 & w4_155;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1120_start: Boolean;
  signal convolution3D_CP_1120_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_576_inst_req_0 : boolean;
  signal type_cast_1234_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_538_inst_ack_0 : boolean;
  signal type_cast_530_inst_req_0 : boolean;
  signal type_cast_617_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_538_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_613_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_576_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_576_inst_req_1 : boolean;
  signal type_cast_630_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_588_inst_ack_1 : boolean;
  signal type_cast_567_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_613_inst_ack_1 : boolean;
  signal type_cast_630_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_563_inst_ack_1 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_588_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_551_inst_ack_1 : boolean;
  signal type_cast_530_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_501_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_551_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_551_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_526_inst_req_1 : boolean;
  signal type_cast_630_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_526_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_613_inst_req_1 : boolean;
  signal type_cast_580_inst_ack_0 : boolean;
  signal type_cast_659_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_588_inst_req_1 : boolean;
  signal type_cast_567_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_613_inst_ack_0 : boolean;
  signal type_cast_617_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_588_inst_req_0 : boolean;
  signal type_cast_530_inst_ack_0 : boolean;
  signal type_cast_617_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_551_inst_ack_0 : boolean;
  signal type_cast_517_inst_req_1 : boolean;
  signal type_cast_505_inst_ack_1 : boolean;
  signal type_cast_505_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_538_inst_ack_1 : boolean;
  signal type_cast_639_inst_ack_1 : boolean;
  signal type_cast_659_inst_req_0 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal type_cast_505_inst_req_1 : boolean;
  signal type_cast_643_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_526_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_538_inst_req_1 : boolean;
  signal type_cast_517_inst_ack_0 : boolean;
  signal type_cast_1265_inst_req_1 : boolean;
  signal type_cast_659_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_576_inst_ack_0 : boolean;
  signal type_cast_505_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_501_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_626_inst_ack_1 : boolean;
  signal type_cast_659_inst_req_1 : boolean;
  signal type_cast_643_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_626_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_563_inst_req_1 : boolean;
  signal type_cast_1301_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_526_inst_req_0 : boolean;
  signal type_cast_1234_inst_req_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_555_inst_req_0 : boolean;
  signal type_cast_555_inst_ack_0 : boolean;
  signal type_cast_630_inst_req_0 : boolean;
  signal type_cast_580_inst_req_1 : boolean;
  signal type_cast_555_inst_req_1 : boolean;
  signal type_cast_530_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_req_0 : boolean;
  signal type_cast_580_inst_req_0 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal type_cast_605_inst_req_0 : boolean;
  signal type_cast_639_inst_req_0 : boolean;
  signal type_cast_605_inst_ack_0 : boolean;
  signal type_cast_555_inst_ack_1 : boolean;
  signal type_cast_639_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_513_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_513_inst_req_0 : boolean;
  signal type_cast_617_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_ack_0 : boolean;
  signal type_cast_1265_inst_req_0 : boolean;
  signal type_cast_687_inst_req_1 : boolean;
  signal type_cast_687_inst_ack_1 : boolean;
  signal type_cast_703_inst_ack_1 : boolean;
  signal type_cast_703_inst_req_1 : boolean;
  signal type_cast_542_inst_ack_1 : boolean;
  signal type_cast_639_inst_req_1 : boolean;
  signal type_cast_687_inst_req_0 : boolean;
  signal type_cast_687_inst_ack_0 : boolean;
  signal type_cast_517_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_626_inst_ack_0 : boolean;
  signal type_cast_567_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_626_inst_req_0 : boolean;
  signal type_cast_712_inst_req_0 : boolean;
  signal type_cast_712_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_req_0 : boolean;
  signal type_cast_542_inst_req_1 : boolean;
  signal type_cast_1265_inst_ack_0 : boolean;
  signal type_cast_567_inst_req_1 : boolean;
  signal if_stmt_667_branch_ack_1 : boolean;
  signal type_cast_592_inst_ack_1 : boolean;
  signal if_stmt_667_branch_ack_0 : boolean;
  signal type_cast_703_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_req_1 : boolean;
  signal type_cast_703_inst_ack_0 : boolean;
  signal type_cast_712_inst_req_1 : boolean;
  signal type_cast_712_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1230_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1230_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_ack_1 : boolean;
  signal if_stmt_667_branch_req_0 : boolean;
  signal type_cast_1301_inst_req_0 : boolean;
  signal type_cast_580_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_563_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_563_inst_req_0 : boolean;
  signal type_cast_1234_inst_req_1 : boolean;
  signal type_cast_542_inst_ack_0 : boolean;
  signal type_cast_542_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_513_inst_ack_1 : boolean;
  signal type_cast_605_inst_ack_1 : boolean;
  signal type_cast_592_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_513_inst_req_1 : boolean;
  signal type_cast_1627_inst_ack_1 : boolean;
  signal type_cast_1234_inst_ack_1 : boolean;
  signal array_obj_ref_1226_index_offset_req_1 : boolean;
  signal type_cast_517_inst_ack_1 : boolean;
  signal array_obj_ref_1226_index_offset_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_ack_1 : boolean;
  signal type_cast_1265_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1243_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1243_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_ack_1 : boolean;
  signal type_cast_1319_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1243_inst_req_1 : boolean;
  signal addr_of_1227_final_reg_req_0 : boolean;
  signal type_cast_442_inst_req_0 : boolean;
  signal type_cast_442_inst_ack_0 : boolean;
  signal type_cast_442_inst_req_1 : boolean;
  signal type_cast_442_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_451_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_451_inst_ack_0 : boolean;
  signal type_cast_1319_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_451_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_451_inst_ack_1 : boolean;
  signal type_cast_455_inst_req_0 : boolean;
  signal type_cast_455_inst_ack_0 : boolean;
  signal type_cast_455_inst_req_1 : boolean;
  signal type_cast_455_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_463_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_463_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_463_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_463_inst_ack_1 : boolean;
  signal type_cast_605_inst_req_1 : boolean;
  signal type_cast_467_inst_req_0 : boolean;
  signal type_cast_467_inst_ack_0 : boolean;
  signal type_cast_467_inst_req_1 : boolean;
  signal type_cast_467_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_476_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_476_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_476_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_476_inst_ack_1 : boolean;
  signal type_cast_480_inst_req_0 : boolean;
  signal type_cast_480_inst_ack_0 : boolean;
  signal type_cast_480_inst_req_1 : boolean;
  signal type_cast_480_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_488_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_488_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_488_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_488_inst_ack_1 : boolean;
  signal type_cast_492_inst_req_0 : boolean;
  signal type_cast_492_inst_ack_0 : boolean;
  signal type_cast_492_inst_req_1 : boolean;
  signal type_cast_492_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_501_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_501_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_req_1 : boolean;
  signal type_cast_1283_inst_ack_1 : boolean;
  signal type_cast_722_inst_req_0 : boolean;
  signal type_cast_1283_inst_req_1 : boolean;
  signal type_cast_722_inst_ack_0 : boolean;
  signal type_cast_722_inst_req_1 : boolean;
  signal type_cast_722_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_req_0 : boolean;
  signal array_obj_ref_1226_index_offset_ack_0 : boolean;
  signal array_obj_ref_757_index_offset_req_0 : boolean;
  signal type_cast_1283_inst_ack_0 : boolean;
  signal array_obj_ref_757_index_offset_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1230_inst_ack_0 : boolean;
  signal array_obj_ref_757_index_offset_req_1 : boolean;
  signal type_cast_1283_inst_req_0 : boolean;
  signal array_obj_ref_757_index_offset_ack_1 : boolean;
  signal type_cast_1247_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1230_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_ack_1 : boolean;
  signal addr_of_758_final_reg_req_0 : boolean;
  signal addr_of_758_final_reg_ack_0 : boolean;
  signal addr_of_758_final_reg_req_1 : boolean;
  signal addr_of_758_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_761_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_761_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_761_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_761_inst_ack_1 : boolean;
  signal type_cast_1247_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_req_1 : boolean;
  signal type_cast_1247_inst_ack_0 : boolean;
  signal type_cast_1247_inst_req_0 : boolean;
  signal type_cast_1319_inst_ack_1 : boolean;
  signal type_cast_765_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_ack_1 : boolean;
  signal type_cast_765_inst_ack_0 : boolean;
  signal type_cast_1319_inst_req_1 : boolean;
  signal type_cast_765_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_req_1 : boolean;
  signal type_cast_765_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_774_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_774_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_774_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_774_inst_ack_1 : boolean;
  signal type_cast_1337_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1243_inst_ack_1 : boolean;
  signal array_obj_ref_1226_index_offset_req_0 : boolean;
  signal type_cast_778_inst_req_0 : boolean;
  signal type_cast_778_inst_ack_0 : boolean;
  signal type_cast_778_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_ack_0 : boolean;
  signal type_cast_778_inst_ack_1 : boolean;
  signal addr_of_1227_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_ack_0 : boolean;
  signal addr_of_1227_final_reg_req_1 : boolean;
  signal type_cast_1301_inst_ack_1 : boolean;
  signal type_cast_1301_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_ack_1 : boolean;
  signal type_cast_1337_inst_req_0 : boolean;
  signal addr_of_1227_final_reg_ack_0 : boolean;
  signal type_cast_1044_inst_req_0 : boolean;
  signal type_cast_1044_inst_ack_0 : boolean;
  signal type_cast_796_inst_req_0 : boolean;
  signal type_cast_796_inst_ack_0 : boolean;
  signal type_cast_796_inst_req_1 : boolean;
  signal type_cast_796_inst_ack_1 : boolean;
  signal phi_stmt_980_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_ack_1 : boolean;
  signal type_cast_1044_inst_req_1 : boolean;
  signal type_cast_814_inst_req_0 : boolean;
  signal type_cast_814_inst_ack_0 : boolean;
  signal type_cast_942_inst_ack_1 : boolean;
  signal type_cast_814_inst_req_1 : boolean;
  signal phi_stmt_939_req_1 : boolean;
  signal type_cast_814_inst_ack_1 : boolean;
  signal phi_stmt_1624_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_req_1 : boolean;
  signal type_cast_1044_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_ack_1 : boolean;
  signal phi_stmt_1624_req_1 : boolean;
  signal phi_stmt_1041_req_0 : boolean;
  signal type_cast_832_inst_req_0 : boolean;
  signal phi_stmt_1408_req_1 : boolean;
  signal type_cast_832_inst_ack_0 : boolean;
  signal type_cast_832_inst_req_1 : boolean;
  signal type_cast_832_inst_ack_1 : boolean;
  signal type_cast_986_inst_ack_1 : boolean;
  signal phi_stmt_1041_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_ack_1 : boolean;
  signal type_cast_850_inst_req_0 : boolean;
  signal type_cast_850_inst_ack_0 : boolean;
  signal type_cast_850_inst_req_1 : boolean;
  signal type_cast_850_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_req_0 : boolean;
  signal phi_stmt_1408_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_ack_1 : boolean;
  signal phi_stmt_987_req_0 : boolean;
  signal phi_stmt_939_req_0 : boolean;
  signal type_cast_868_inst_req_0 : boolean;
  signal type_cast_868_inst_ack_0 : boolean;
  signal type_cast_868_inst_req_1 : boolean;
  signal type_cast_868_inst_ack_1 : boolean;
  signal phi_stmt_980_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_ack_1 : boolean;
  signal type_cast_886_inst_req_0 : boolean;
  signal type_cast_886_inst_ack_0 : boolean;
  signal type_cast_886_inst_req_1 : boolean;
  signal type_cast_886_inst_ack_1 : boolean;
  signal type_cast_1459_inst_req_0 : boolean;
  signal type_cast_1459_inst_ack_0 : boolean;
  signal ptr_deref_894_store_0_req_0 : boolean;
  signal ptr_deref_894_store_0_ack_0 : boolean;
  signal phi_stmt_939_ack_0 : boolean;
  signal ptr_deref_894_store_0_req_1 : boolean;
  signal ptr_deref_894_store_0_ack_1 : boolean;
  signal type_cast_1220_inst_req_0 : boolean;
  signal if_stmt_908_branch_req_0 : boolean;
  signal if_stmt_908_branch_ack_1 : boolean;
  signal if_stmt_908_branch_ack_0 : boolean;
  signal type_cast_1220_inst_ack_0 : boolean;
  signal type_cast_1517_inst_req_0 : boolean;
  signal type_cast_1517_inst_ack_0 : boolean;
  signal if_stmt_959_branch_req_0 : boolean;
  signal if_stmt_959_branch_ack_1 : boolean;
  signal if_stmt_959_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1008_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1008_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1008_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1008_inst_ack_1 : boolean;
  signal type_cast_1012_inst_req_0 : boolean;
  signal type_cast_1012_inst_ack_0 : boolean;
  signal type_cast_1012_inst_req_1 : boolean;
  signal type_cast_1012_inst_ack_1 : boolean;
  signal type_cast_1027_inst_req_0 : boolean;
  signal phi_stmt_1214_req_0 : boolean;
  signal type_cast_1027_inst_ack_0 : boolean;
  signal type_cast_1027_inst_req_1 : boolean;
  signal type_cast_1027_inst_ack_1 : boolean;
  signal type_cast_986_inst_req_0 : boolean;
  signal type_cast_1459_inst_req_1 : boolean;
  signal type_cast_942_inst_req_0 : boolean;
  signal if_stmt_1034_branch_req_0 : boolean;
  signal if_stmt_1034_branch_ack_1 : boolean;
  signal if_stmt_1034_branch_ack_0 : boolean;
  signal array_obj_ref_1073_index_offset_req_0 : boolean;
  signal array_obj_ref_1073_index_offset_ack_0 : boolean;
  signal array_obj_ref_1073_index_offset_req_1 : boolean;
  signal array_obj_ref_1073_index_offset_ack_1 : boolean;
  signal addr_of_1074_final_reg_req_0 : boolean;
  signal addr_of_1074_final_reg_ack_0 : boolean;
  signal addr_of_1074_final_reg_req_1 : boolean;
  signal addr_of_1074_final_reg_ack_1 : boolean;
  signal ptr_deref_1077_store_0_req_0 : boolean;
  signal ptr_deref_1077_store_0_ack_0 : boolean;
  signal ptr_deref_1077_store_0_req_1 : boolean;
  signal ptr_deref_1077_store_0_ack_1 : boolean;
  signal type_cast_1084_inst_req_0 : boolean;
  signal type_cast_1084_inst_ack_0 : boolean;
  signal type_cast_1084_inst_req_1 : boolean;
  signal type_cast_1084_inst_ack_1 : boolean;
  signal type_cast_1088_inst_req_0 : boolean;
  signal type_cast_1088_inst_ack_0 : boolean;
  signal type_cast_1088_inst_req_1 : boolean;
  signal type_cast_1088_inst_ack_1 : boolean;
  signal type_cast_1092_inst_req_0 : boolean;
  signal type_cast_1092_inst_ack_0 : boolean;
  signal type_cast_1092_inst_req_1 : boolean;
  signal type_cast_1092_inst_ack_1 : boolean;
  signal type_cast_1096_inst_req_0 : boolean;
  signal type_cast_1096_inst_ack_0 : boolean;
  signal type_cast_1096_inst_req_1 : boolean;
  signal type_cast_1096_inst_ack_1 : boolean;
  signal if_stmt_1134_branch_req_0 : boolean;
  signal if_stmt_1134_branch_ack_1 : boolean;
  signal if_stmt_1134_branch_ack_0 : boolean;
  signal type_cast_1155_inst_req_0 : boolean;
  signal type_cast_1155_inst_ack_0 : boolean;
  signal type_cast_1155_inst_req_1 : boolean;
  signal type_cast_1155_inst_ack_1 : boolean;
  signal type_cast_1159_inst_req_0 : boolean;
  signal type_cast_1159_inst_ack_0 : boolean;
  signal type_cast_1159_inst_req_1 : boolean;
  signal type_cast_1159_inst_ack_1 : boolean;
  signal type_cast_1168_inst_req_0 : boolean;
  signal type_cast_1168_inst_ack_0 : boolean;
  signal type_cast_1168_inst_req_1 : boolean;
  signal type_cast_1168_inst_ack_1 : boolean;
  signal type_cast_1177_inst_req_0 : boolean;
  signal type_cast_1177_inst_ack_0 : boolean;
  signal type_cast_1177_inst_req_1 : boolean;
  signal type_cast_1177_inst_ack_1 : boolean;
  signal type_cast_1186_inst_req_0 : boolean;
  signal type_cast_1186_inst_ack_0 : boolean;
  signal type_cast_1186_inst_req_1 : boolean;
  signal type_cast_1186_inst_ack_1 : boolean;
  signal type_cast_1191_inst_req_0 : boolean;
  signal type_cast_1191_inst_ack_0 : boolean;
  signal type_cast_1191_inst_req_1 : boolean;
  signal type_cast_1191_inst_ack_1 : boolean;
  signal type_cast_1337_inst_req_1 : boolean;
  signal type_cast_1337_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_ack_1 : boolean;
  signal type_cast_1355_inst_req_0 : boolean;
  signal type_cast_1355_inst_ack_0 : boolean;
  signal type_cast_1355_inst_req_1 : boolean;
  signal type_cast_1355_inst_ack_1 : boolean;
  signal ptr_deref_1363_store_0_req_0 : boolean;
  signal ptr_deref_1363_store_0_ack_0 : boolean;
  signal ptr_deref_1363_store_0_req_1 : boolean;
  signal ptr_deref_1363_store_0_ack_1 : boolean;
  signal if_stmt_1377_branch_req_0 : boolean;
  signal if_stmt_1377_branch_ack_1 : boolean;
  signal if_stmt_1377_branch_ack_0 : boolean;
  signal if_stmt_1428_branch_req_0 : boolean;
  signal if_stmt_1428_branch_ack_1 : boolean;
  signal if_stmt_1428_branch_ack_0 : boolean;
  signal type_cast_1443_inst_req_0 : boolean;
  signal type_cast_1443_inst_ack_0 : boolean;
  signal type_cast_1443_inst_req_1 : boolean;
  signal type_cast_1443_inst_ack_1 : boolean;
  signal type_cast_1627_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1481_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1481_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1481_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1481_inst_ack_1 : boolean;
  signal type_cast_1466_inst_ack_0 : boolean;
  signal type_cast_1485_inst_req_0 : boolean;
  signal phi_stmt_1408_req_0 : boolean;
  signal type_cast_1485_inst_ack_0 : boolean;
  signal type_cast_1485_inst_req_1 : boolean;
  signal type_cast_1411_inst_ack_1 : boolean;
  signal type_cast_1485_inst_ack_1 : boolean;
  signal type_cast_1627_inst_ack_0 : boolean;
  signal type_cast_1500_inst_req_0 : boolean;
  signal type_cast_1411_inst_req_1 : boolean;
  signal type_cast_1500_inst_ack_0 : boolean;
  signal type_cast_1500_inst_req_1 : boolean;
  signal type_cast_1500_inst_ack_1 : boolean;
  signal type_cast_1627_inst_req_0 : boolean;
  signal type_cast_942_inst_req_1 : boolean;
  signal if_stmt_1507_branch_req_0 : boolean;
  signal type_cast_1411_inst_ack_0 : boolean;
  signal type_cast_1411_inst_req_0 : boolean;
  signal if_stmt_1507_branch_ack_1 : boolean;
  signal if_stmt_1507_branch_ack_0 : boolean;
  signal type_cast_1466_inst_req_0 : boolean;
  signal type_cast_986_inst_req_1 : boolean;
  signal array_obj_ref_1546_index_offset_req_0 : boolean;
  signal array_obj_ref_1546_index_offset_ack_0 : boolean;
  signal array_obj_ref_1546_index_offset_req_1 : boolean;
  signal array_obj_ref_1546_index_offset_ack_1 : boolean;
  signal addr_of_1547_final_reg_req_0 : boolean;
  signal addr_of_1547_final_reg_ack_0 : boolean;
  signal addr_of_1547_final_reg_req_1 : boolean;
  signal addr_of_1547_final_reg_ack_1 : boolean;
  signal phi_stmt_1460_req_0 : boolean;
  signal ptr_deref_1550_store_0_req_0 : boolean;
  signal phi_stmt_987_ack_0 : boolean;
  signal ptr_deref_1550_store_0_ack_0 : boolean;
  signal type_cast_942_inst_ack_0 : boolean;
  signal type_cast_986_inst_ack_0 : boolean;
  signal ptr_deref_1550_store_0_req_1 : boolean;
  signal phi_stmt_980_ack_0 : boolean;
  signal ptr_deref_1550_store_0_ack_1 : boolean;
  signal phi_stmt_1453_req_0 : boolean;
  signal call_stmt_1557_call_req_0 : boolean;
  signal call_stmt_1557_call_ack_0 : boolean;
  signal call_stmt_1557_call_req_1 : boolean;
  signal call_stmt_1557_call_ack_1 : boolean;
  signal phi_stmt_1514_ack_0 : boolean;
  signal phi_stmt_1453_req_1 : boolean;
  signal WPIPE_num_out_pipe_1569_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1569_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1569_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1569_inst_ack_1 : boolean;
  signal phi_stmt_1514_req_0 : boolean;
  signal phi_stmt_987_req_1 : boolean;
  signal type_cast_993_inst_ack_1 : boolean;
  signal type_cast_1459_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1572_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1572_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1572_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1572_inst_ack_1 : boolean;
  signal type_cast_1466_inst_req_1 : boolean;
  signal type_cast_1517_inst_ack_1 : boolean;
  signal type_cast_993_inst_req_1 : boolean;
  signal type_cast_1517_inst_req_1 : boolean;
  signal type_cast_993_inst_ack_0 : boolean;
  signal phi_stmt_1460_ack_0 : boolean;
  signal type_cast_1596_inst_req_0 : boolean;
  signal phi_stmt_1214_ack_0 : boolean;
  signal type_cast_1596_inst_ack_0 : boolean;
  signal phi_stmt_1453_ack_0 : boolean;
  signal type_cast_1596_inst_req_1 : boolean;
  signal type_cast_1596_inst_ack_1 : boolean;
  signal type_cast_993_inst_req_0 : boolean;
  signal type_cast_1606_inst_req_0 : boolean;
  signal type_cast_1606_inst_ack_0 : boolean;
  signal type_cast_1606_inst_req_1 : boolean;
  signal phi_stmt_1214_req_1 : boolean;
  signal type_cast_1606_inst_ack_1 : boolean;
  signal phi_stmt_1460_req_1 : boolean;
  signal type_cast_1615_inst_req_0 : boolean;
  signal type_cast_1220_inst_ack_1 : boolean;
  signal type_cast_1615_inst_ack_0 : boolean;
  signal type_cast_1466_inst_ack_1 : boolean;
  signal type_cast_1615_inst_req_1 : boolean;
  signal type_cast_1220_inst_req_1 : boolean;
  signal type_cast_1615_inst_ack_1 : boolean;
  signal type_cast_1644_inst_req_0 : boolean;
  signal type_cast_1644_inst_ack_0 : boolean;
  signal type_cast_1644_inst_req_1 : boolean;
  signal type_cast_1644_inst_ack_1 : boolean;
  signal type_cast_1648_inst_req_0 : boolean;
  signal type_cast_1648_inst_ack_0 : boolean;
  signal type_cast_1648_inst_req_1 : boolean;
  signal type_cast_1648_inst_ack_1 : boolean;
  signal call_stmt_1652_call_req_0 : boolean;
  signal call_stmt_1652_call_ack_0 : boolean;
  signal call_stmt_1652_call_req_1 : boolean;
  signal call_stmt_1652_call_ack_1 : boolean;
  signal call_stmt_1659_call_req_0 : boolean;
  signal call_stmt_1659_call_ack_0 : boolean;
  signal call_stmt_1659_call_req_1 : boolean;
  signal call_stmt_1659_call_ack_1 : boolean;
  signal if_stmt_1671_branch_req_0 : boolean;
  signal if_stmt_1671_branch_ack_1 : boolean;
  signal if_stmt_1671_branch_ack_0 : boolean;
  signal type_cast_1681_inst_req_0 : boolean;
  signal type_cast_1681_inst_ack_0 : boolean;
  signal type_cast_1681_inst_req_1 : boolean;
  signal type_cast_1681_inst_ack_1 : boolean;
  signal call_stmt_1685_call_req_0 : boolean;
  signal call_stmt_1685_call_ack_0 : boolean;
  signal call_stmt_1685_call_req_1 : boolean;
  signal call_stmt_1685_call_ack_1 : boolean;
  signal type_cast_1689_inst_req_0 : boolean;
  signal type_cast_1689_inst_ack_0 : boolean;
  signal type_cast_1689_inst_req_1 : boolean;
  signal type_cast_1689_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1696_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1696_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1696_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1696_inst_ack_1 : boolean;
  signal phi_stmt_745_req_0 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal type_cast_751_inst_req_1 : boolean;
  signal type_cast_751_inst_ack_1 : boolean;
  signal phi_stmt_745_req_1 : boolean;
  signal phi_stmt_745_ack_0 : boolean;
  signal phi_stmt_1624_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1120_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1120: Block -- control-path 
    signal convolution3D_CP_1120_elements: BooleanArray(333 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1120_elements(0) <= convolution3D_CP_1120_start;
    convolution3D_CP_1120_symbol <= convolution3D_CP_1120_elements(265);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_436/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/branch_block_stmt_436__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Update/cr
      -- 
    cr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_630_inst_req_1); -- 
    cr_1451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_530_inst_req_1); -- 
    cr_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_617_inst_req_1); -- 
    cr_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_517_inst_req_1); -- 
    cr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_505_inst_req_1); -- 
    cr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_659_inst_req_1); -- 
    cr_1703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_643_inst_req_1); -- 
    cr_1563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_580_inst_req_1); -- 
    cr_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_555_inst_req_1); -- 
    cr_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_639_inst_req_1); -- 
    cr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_542_inst_req_1); -- 
    cr_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_567_inst_req_1); -- 
    cr_1591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_592_inst_req_1); -- 
    rr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => RPIPE_maxpool_input_pipe_438_inst_req_0); -- 
    cr_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_442_inst_req_1); -- 
    cr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_455_inst_req_1); -- 
    cr_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_605_inst_req_1); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_467_inst_req_1); -- 
    cr_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_480_inst_req_1); -- 
    cr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_492_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_update_start_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Update/cr
      -- 
    ra_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_438_inst_ack_0, ack => convolution3D_CP_1120_elements(1)); -- 
    cr_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(1), ack => RPIPE_maxpool_input_pipe_438_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_438_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Sample/rr
      -- 
    ca_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_438_inst_ack_1, ack => convolution3D_CP_1120_elements(2)); -- 
    rr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => type_cast_442_inst_req_0); -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => RPIPE_maxpool_input_pipe_451_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Sample/ra
      -- 
    ra_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_442_inst_ack_0, ack => convolution3D_CP_1120_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_442_Update/ca
      -- 
    ca_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_442_inst_ack_1, ack => convolution3D_CP_1120_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_update_start_
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Update/cr
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_451_inst_ack_0, ack => convolution3D_CP_1120_elements(5)); -- 
    cr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(5), ack => RPIPE_maxpool_input_pipe_451_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_451_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Sample/rr
      -- 
    ca_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_451_inst_ack_1, ack => convolution3D_CP_1120_elements(6)); -- 
    rr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => type_cast_455_inst_req_0); -- 
    rr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => RPIPE_maxpool_input_pipe_463_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Sample/ra
      -- 
    ra_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_455_inst_ack_0, ack => convolution3D_CP_1120_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_455_Update/ca
      -- 
    ca_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_455_inst_ack_1, ack => convolution3D_CP_1120_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_update_start_
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Update/cr
      -- 
    ra_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_463_inst_ack_0, ack => convolution3D_CP_1120_elements(9)); -- 
    cr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(9), ack => RPIPE_maxpool_input_pipe_463_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_463_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Sample/rr
      -- 
    ca_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_463_inst_ack_1, ack => convolution3D_CP_1120_elements(10)); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(10), ack => type_cast_467_inst_req_0); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(10), ack => RPIPE_maxpool_input_pipe_476_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Sample/ra
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_467_inst_ack_0, ack => convolution3D_CP_1120_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_467_Update/ca
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_467_inst_ack_1, ack => convolution3D_CP_1120_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_update_start_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Update/cr
      -- 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_476_inst_ack_0, ack => convolution3D_CP_1120_elements(13)); -- 
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(13), ack => RPIPE_maxpool_input_pipe_476_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_476_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Sample/rr
      -- 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_476_inst_ack_1, ack => convolution3D_CP_1120_elements(14)); -- 
    rr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(14), ack => type_cast_480_inst_req_0); -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(14), ack => RPIPE_maxpool_input_pipe_488_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Sample/ra
      -- 
    ra_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_0, ack => convolution3D_CP_1120_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_480_Update/ca
      -- 
    ca_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_1, ack => convolution3D_CP_1120_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_update_start_
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Update/cr
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_488_inst_ack_0, ack => convolution3D_CP_1120_elements(17)); -- 
    cr_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(17), ack => RPIPE_maxpool_input_pipe_488_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_488_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Sample/rr
      -- 
    ca_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_488_inst_ack_1, ack => convolution3D_CP_1120_elements(18)); -- 
    rr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(18), ack => type_cast_492_inst_req_0); -- 
    rr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(18), ack => RPIPE_maxpool_input_pipe_501_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Sample/ra
      -- 
    ra_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_0, ack => convolution3D_CP_1120_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_492_Update/ca
      -- 
    ca_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_1, ack => convolution3D_CP_1120_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_update_start_
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Sample/ra
      -- 
    ra_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_501_inst_ack_0, ack => convolution3D_CP_1120_elements(21)); -- 
    cr_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(21), ack => RPIPE_maxpool_input_pipe_501_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_501_update_completed_
      -- 
    ca_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_501_inst_ack_1, ack => convolution3D_CP_1120_elements(22)); -- 
    rr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(22), ack => type_cast_505_inst_req_0); -- 
    rr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(22), ack => RPIPE_maxpool_input_pipe_513_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Sample/$exit
      -- 
    ra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_505_inst_ack_0, ack => convolution3D_CP_1120_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_505_Update/$exit
      -- 
    ca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_505_inst_ack_1, ack => convolution3D_CP_1120_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_update_start_
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Update/cr
      -- 
    ra_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_513_inst_ack_0, ack => convolution3D_CP_1120_elements(25)); -- 
    cr_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(25), ack => RPIPE_maxpool_input_pipe_513_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_513_Update/$exit
      -- 
    ca_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_513_inst_ack_1, ack => convolution3D_CP_1120_elements(26)); -- 
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(26), ack => type_cast_517_inst_req_0); -- 
    rr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(26), ack => RPIPE_maxpool_input_pipe_526_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_sample_completed_
      -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_517_inst_ack_0, ack => convolution3D_CP_1120_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_517_Update/ca
      -- 
    ca_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_517_inst_ack_1, ack => convolution3D_CP_1120_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_update_start_
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_sample_completed_
      -- 
    ra_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_526_inst_ack_0, ack => convolution3D_CP_1120_elements(29)); -- 
    cr_1437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(29), ack => RPIPE_maxpool_input_pipe_526_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_526_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_sample_start_
      -- 
    ca_1438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_526_inst_ack_1, ack => convolution3D_CP_1120_elements(30)); -- 
    rr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(30), ack => type_cast_530_inst_req_0); -- 
    rr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(30), ack => RPIPE_maxpool_input_pipe_538_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_sample_completed_
      -- 
    ra_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_530_inst_ack_0, ack => convolution3D_CP_1120_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_530_Update/ca
      -- 
    ca_1452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_530_inst_ack_1, ack => convolution3D_CP_1120_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_update_start_
      -- 
    ra_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_538_inst_ack_0, ack => convolution3D_CP_1120_elements(33)); -- 
    cr_1465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(33), ack => RPIPE_maxpool_input_pipe_538_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_538_update_completed_
      -- 
    ca_1466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_538_inst_ack_1, ack => convolution3D_CP_1120_elements(34)); -- 
    rr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(34), ack => type_cast_542_inst_req_0); -- 
    rr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(34), ack => RPIPE_maxpool_input_pipe_551_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Sample/$exit
      -- 
    ra_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_0, ack => convolution3D_CP_1120_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_542_Update/$exit
      -- 
    ca_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_1, ack => convolution3D_CP_1120_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_update_start_
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_sample_completed_
      -- 
    ra_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_551_inst_ack_0, ack => convolution3D_CP_1120_elements(37)); -- 
    cr_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(37), ack => RPIPE_maxpool_input_pipe_551_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_551_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Sample/$entry
      -- 
    ca_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_551_inst_ack_1, ack => convolution3D_CP_1120_elements(38)); -- 
    rr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(38), ack => type_cast_555_inst_req_0); -- 
    rr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(38), ack => RPIPE_maxpool_input_pipe_563_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Sample/ra
      -- 
    ra_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_555_inst_ack_0, ack => convolution3D_CP_1120_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_555_Update/ca
      -- 
    ca_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_555_inst_ack_1, ack => convolution3D_CP_1120_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_update_start_
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Sample/$exit
      -- 
    ra_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_563_inst_ack_0, ack => convolution3D_CP_1120_elements(41)); -- 
    cr_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(41), ack => RPIPE_maxpool_input_pipe_563_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_563_update_completed_
      -- 
    ca_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_563_inst_ack_1, ack => convolution3D_CP_1120_elements(42)); -- 
    rr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => type_cast_567_inst_req_0); -- 
    rr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => RPIPE_maxpool_input_pipe_576_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Sample/ra
      -- 
    ra_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_567_inst_ack_0, ack => convolution3D_CP_1120_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_567_Update/$exit
      -- 
    ca_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_567_inst_ack_1, ack => convolution3D_CP_1120_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Update/cr
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_update_start_
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Sample/ra
      -- 
    ra_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_576_inst_ack_0, ack => convolution3D_CP_1120_elements(45)); -- 
    cr_1549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(45), ack => RPIPE_maxpool_input_pipe_576_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_576_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_sample_start_
      -- 
    ca_1550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_576_inst_ack_1, ack => convolution3D_CP_1120_elements(46)); -- 
    rr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(46), ack => type_cast_580_inst_req_0); -- 
    rr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(46), ack => RPIPE_maxpool_input_pipe_588_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_sample_completed_
      -- 
    ra_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_580_inst_ack_0, ack => convolution3D_CP_1120_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_580_Update/ca
      -- 
    ca_1564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_580_inst_ack_1, ack => convolution3D_CP_1120_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_update_start_
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_sample_completed_
      -- 
    ra_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_588_inst_ack_0, ack => convolution3D_CP_1120_elements(49)); -- 
    cr_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(49), ack => RPIPE_maxpool_input_pipe_588_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_588_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_sample_start_
      -- 
    ca_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_588_inst_ack_1, ack => convolution3D_CP_1120_elements(50)); -- 
    rr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => type_cast_592_inst_req_0); -- 
    rr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => RPIPE_maxpool_input_pipe_601_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Sample/ra
      -- 
    ra_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => convolution3D_CP_1120_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_592_Update/ca
      -- 
    ca_1592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_1, ack => convolution3D_CP_1120_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_update_start_
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_sample_completed_
      -- 
    ra_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_601_inst_ack_0, ack => convolution3D_CP_1120_elements(53)); -- 
    cr_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(53), ack => RPIPE_maxpool_input_pipe_601_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_601_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_sample_start_
      -- 
    ca_1606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_601_inst_ack_1, ack => convolution3D_CP_1120_elements(54)); -- 
    rr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(54), ack => type_cast_605_inst_req_0); -- 
    rr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(54), ack => RPIPE_maxpool_input_pipe_613_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Sample/ra
      -- 
    ra_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_605_inst_ack_0, ack => convolution3D_CP_1120_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_605_Update/ca
      -- 
    ca_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_605_inst_ack_1, ack => convolution3D_CP_1120_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_update_start_
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_sample_completed_
      -- 
    ra_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_613_inst_ack_0, ack => convolution3D_CP_1120_elements(57)); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(57), ack => RPIPE_maxpool_input_pipe_613_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_613_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Sample/$entry
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_613_inst_ack_1, ack => convolution3D_CP_1120_elements(58)); -- 
    rr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(58), ack => type_cast_617_inst_req_0); -- 
    rr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(58), ack => RPIPE_maxpool_input_pipe_626_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Sample/ra
      -- 
    ra_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_617_inst_ack_0, ack => convolution3D_CP_1120_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_617_Update/$exit
      -- 
    ca_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_617_inst_ack_1, ack => convolution3D_CP_1120_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_update_start_
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Update/cr
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Sample/$exit
      -- 
    ra_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_626_inst_ack_0, ack => convolution3D_CP_1120_elements(61)); -- 
    cr_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(61), ack => RPIPE_maxpool_input_pipe_626_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/RPIPE_maxpool_input_pipe_626_update_completed_
      -- 
    ca_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_626_inst_ack_1, ack => convolution3D_CP_1120_elements(62)); -- 
    rr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(62), ack => type_cast_630_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Sample/$exit
      -- 
    ra_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_630_inst_ack_0, ack => convolution3D_CP_1120_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_630_Update/$exit
      -- 
    ca_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_630_inst_ack_1, ack => convolution3D_CP_1120_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Sample/rr
      -- 
    rr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(65), ack => type_cast_639_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(12) & convolution3D_CP_1120_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Sample/ra
      -- 
    ra_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_0, ack => convolution3D_CP_1120_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_639_Update/$exit
      -- 
    ca_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_1, ack => convolution3D_CP_1120_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_sample_start_
      -- 
    rr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(68), ack => type_cast_643_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(20) & convolution3D_CP_1120_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_sample_completed_
      -- 
    ra_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => convolution3D_CP_1120_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_643_Update/ca
      -- 
    ca_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_1, ack => convolution3D_CP_1120_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Sample/$entry
      -- 
    rr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(71), ack => type_cast_659_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(4) & convolution3D_CP_1120_elements(8) & convolution3D_CP_1120_elements(67) & convolution3D_CP_1120_elements(70);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Sample/$exit
      -- 
    ra_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_0, ack => convolution3D_CP_1120_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/type_cast_659_update_completed_
      -- 
    ca_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_1, ack => convolution3D_CP_1120_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_667_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_667_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_667_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_667_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_667_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_667_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_436/R_cmp321_668_place
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666__exit__
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_667__entry__
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_666/$exit
      -- 
    branch_req_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(74), ack => if_stmt_667_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(28) & convolution3D_CP_1120_elements(32) & convolution3D_CP_1120_elements(36) & convolution3D_CP_1120_elements(40) & convolution3D_CP_1120_elements(44) & convolution3D_CP_1120_elements(48) & convolution3D_CP_1120_elements(52) & convolution3D_CP_1120_elements(56) & convolution3D_CP_1120_elements(60) & convolution3D_CP_1120_elements(64) & convolution3D_CP_1120_elements(73);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/if_stmt_667_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_436/if_stmt_667_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/entry_bbx_xnph323
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_673__exit__
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742__entry__
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/entry_bbx_xnph323_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/entry_bbx_xnph323_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_673_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_673_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_673_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_673_PhiAck/dummy
      -- 
    if_choice_transition_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_667_branch_ack_1, ack => convolution3D_CP_1120_elements(75)); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_687_inst_req_1); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_703_inst_req_1); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_687_inst_req_0); -- 
    rr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_712_inst_req_0); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_703_inst_req_0); -- 
    cr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_712_inst_req_1); -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_722_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	272 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_436/if_stmt_667_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_436/if_stmt_667_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_939/$entry
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$entry
      -- 
    else_choice_transition_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_667_branch_ack_0, ack => convolution3D_CP_1120_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_sample_completed_
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_0, ack => convolution3D_CP_1120_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_687_Update/$exit
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_1, ack => convolution3D_CP_1120_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Sample/ra
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_703_inst_ack_0, ack => convolution3D_CP_1120_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_703_update_completed_
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_703_inst_ack_1, ack => convolution3D_CP_1120_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Sample/ra
      -- 
    ra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_0, ack => convolution3D_CP_1120_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_712_Update/ca
      -- 
    ca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_1, ack => convolution3D_CP_1120_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Sample/rr
      -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(83), ack => type_cast_722_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(80) & convolution3D_CP_1120_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Sample/ra
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_0, ack => convolution3D_CP_1120_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/type_cast_722_Update/ca
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_1, ack => convolution3D_CP_1120_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	266 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742/$exit
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_678_to_assign_stmt_742__exit__
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_745/$entry
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(78) & convolution3D_CP_1120_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	271 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Sample/ack
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_757_index_offset_ack_0, ack => convolution3D_CP_1120_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	271 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_request/req
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_757_index_offset_ack_1, ack => convolution3D_CP_1120_elements(88)); -- 
    req_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(88), ack => addr_of_758_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_request/ack
      -- 
    ack_1840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_758_final_reg_ack_0, ack => convolution3D_CP_1120_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	271 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_word_addrgen/root_register_ack
      -- 
    ack_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_758_final_reg_ack_1, ack => convolution3D_CP_1120_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	271 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_update_start_
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Update/cr
      -- 
    ra_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_761_inst_ack_0, ack => convolution3D_CP_1120_elements(91)); -- 
    cr_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(91), ack => RPIPE_maxpool_input_pipe_761_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Sample/rr
      -- 
    ca_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_761_inst_ack_1, ack => convolution3D_CP_1120_elements(92)); -- 
    rr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(92), ack => type_cast_765_inst_req_0); -- 
    rr_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(92), ack => RPIPE_maxpool_input_pipe_774_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Sample/ra
      -- 
    ra_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_765_inst_ack_0, ack => convolution3D_CP_1120_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	271 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Update/ca
      -- 
    ca_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_765_inst_ack_1, ack => convolution3D_CP_1120_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_update_start_
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Update/cr
      -- 
    ra_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_774_inst_ack_0, ack => convolution3D_CP_1120_elements(95)); -- 
    cr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(95), ack => RPIPE_maxpool_input_pipe_774_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_774_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Sample/rr
      -- 
    ca_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_774_inst_ack_1, ack => convolution3D_CP_1120_elements(96)); -- 
    rr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(96), ack => type_cast_778_inst_req_0); -- 
    rr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(96), ack => RPIPE_maxpool_input_pipe_792_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Sample/ra
      -- 
    ra_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_0, ack => convolution3D_CP_1120_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	271 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Update/ca
      -- 
    ca_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_1, ack => convolution3D_CP_1120_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_update_start_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Update/cr
      -- 
    ra_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_792_inst_ack_0, ack => convolution3D_CP_1120_elements(99)); -- 
    cr_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(99), ack => RPIPE_maxpool_input_pipe_792_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_792_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Sample/rr
      -- 
    ca_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_792_inst_ack_1, ack => convolution3D_CP_1120_elements(100)); -- 
    rr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(100), ack => type_cast_796_inst_req_0); -- 
    rr_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(100), ack => RPIPE_maxpool_input_pipe_810_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Sample/ra
      -- 
    ra_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_796_inst_ack_0, ack => convolution3D_CP_1120_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	271 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Update/ca
      -- 
    ca_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_796_inst_ack_1, ack => convolution3D_CP_1120_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_update_start_
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Update/cr
      -- 
    ra_1938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_810_inst_ack_0, ack => convolution3D_CP_1120_elements(103)); -- 
    cr_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(103), ack => RPIPE_maxpool_input_pipe_810_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_810_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Sample/rr
      -- 
    ca_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_810_inst_ack_1, ack => convolution3D_CP_1120_elements(104)); -- 
    rr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(104), ack => type_cast_814_inst_req_0); -- 
    rr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(104), ack => RPIPE_maxpool_input_pipe_828_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Sample/ra
      -- 
    ra_1952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_0, ack => convolution3D_CP_1120_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	271 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Update/ca
      -- 
    ca_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_1, ack => convolution3D_CP_1120_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_update_start_
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Update/cr
      -- 
    ra_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_828_inst_ack_0, ack => convolution3D_CP_1120_elements(107)); -- 
    cr_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(107), ack => RPIPE_maxpool_input_pipe_828_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_828_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Sample/rr
      -- 
    ca_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_828_inst_ack_1, ack => convolution3D_CP_1120_elements(108)); -- 
    rr_1979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(108), ack => type_cast_832_inst_req_0); -- 
    rr_1993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(108), ack => RPIPE_maxpool_input_pipe_846_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Sample/ra
      -- 
    ra_1980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_0, ack => convolution3D_CP_1120_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	271 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Update/ca
      -- 
    ca_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_1, ack => convolution3D_CP_1120_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_update_start_
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Update/cr
      -- 
    ra_1994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_846_inst_ack_0, ack => convolution3D_CP_1120_elements(111)); -- 
    cr_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(111), ack => RPIPE_maxpool_input_pipe_846_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_846_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Sample/rr
      -- 
    ca_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_846_inst_ack_1, ack => convolution3D_CP_1120_elements(112)); -- 
    rr_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(112), ack => type_cast_850_inst_req_0); -- 
    rr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(112), ack => RPIPE_maxpool_input_pipe_864_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Sample/ra
      -- 
    ra_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_0, ack => convolution3D_CP_1120_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	271 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Update/ca
      -- 
    ca_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_1, ack => convolution3D_CP_1120_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_update_start_
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Update/cr
      -- 
    ra_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_864_inst_ack_0, ack => convolution3D_CP_1120_elements(115)); -- 
    cr_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(115), ack => RPIPE_maxpool_input_pipe_864_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_864_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Sample/rr
      -- 
    ca_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_864_inst_ack_1, ack => convolution3D_CP_1120_elements(116)); -- 
    rr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(116), ack => type_cast_868_inst_req_0); -- 
    rr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(116), ack => RPIPE_maxpool_input_pipe_882_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Sample/ra
      -- 
    ra_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_868_inst_ack_0, ack => convolution3D_CP_1120_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	271 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Update/ca
      -- 
    ca_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_868_inst_ack_1, ack => convolution3D_CP_1120_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_update_start_
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Update/cr
      -- 
    ra_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_882_inst_ack_0, ack => convolution3D_CP_1120_elements(119)); -- 
    cr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(119), ack => RPIPE_maxpool_input_pipe_882_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_882_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Sample/rr
      -- 
    ca_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_882_inst_ack_1, ack => convolution3D_CP_1120_elements(120)); -- 
    rr_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(120), ack => type_cast_886_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Sample/ra
      -- 
    ra_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_886_inst_ack_0, ack => convolution3D_CP_1120_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	271 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Update/ca
      -- 
    ca_2069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_886_inst_ack_1, ack => convolution3D_CP_1120_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/ptr_deref_894_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/ptr_deref_894_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/ptr_deref_894_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/ptr_deref_894_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/word_access_start/word_0/rr
      -- 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(123), ack => ptr_deref_894_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(90) & convolution3D_CP_1120_elements(94) & convolution3D_CP_1120_elements(98) & convolution3D_CP_1120_elements(102) & convolution3D_CP_1120_elements(106) & convolution3D_CP_1120_elements(110) & convolution3D_CP_1120_elements(114) & convolution3D_CP_1120_elements(118) & convolution3D_CP_1120_elements(122);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Sample/word_access_start/word_0/ra
      -- 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_894_store_0_ack_0, ack => convolution3D_CP_1120_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	271 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/word_access_complete/word_0/ca
      -- 
    ca_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_894_store_0_ack_1, ack => convolution3D_CP_1120_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	87 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907__exit__
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_908__entry__
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/$exit
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_908_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_908_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_908_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_908_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_436/R_exitcond32_909_place
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_908_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_908_else_link/$entry
      -- 
    branch_req_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(126), ack => if_stmt_908_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(87) & convolution3D_CP_1120_elements(125);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	273 
    -- CP-element group 127: 	274 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_914__exit__
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_921_to_assign_stmt_936__entry__
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_921_to_assign_stmt_936__exit__
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/if_stmt_908_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/if_stmt_908_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_921_to_assign_stmt_936/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_921_to_assign_stmt_936/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Update/cr
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_914_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_914_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_914_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_914_PhiAck/dummy
      -- 
    if_choice_transition_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_908_branch_ack_1, ack => convolution3D_CP_1120_elements(127)); -- 
    rr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_942_inst_req_0); -- 
    cr_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_942_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	267 
    -- CP-element group 128: 	268 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_436/if_stmt_908_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_436/if_stmt_908_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_908_branch_ack_0, ack => convolution3D_CP_1120_elements(128)); -- 
    rr_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(128), ack => type_cast_751_inst_req_0); -- 
    cr_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(128), ack => type_cast_751_inst_req_1); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	277 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	296 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_436/if_stmt_959_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_436/if_stmt_959_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_436/forx_xend_ifx_xend
      -- 
    if_choice_transition_2157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_959_branch_ack_1, ack => convolution3D_CP_1120_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	277 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	278 
    -- CP-element group 130: 	279 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_965__exit__
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_971_to_assign_stmt_977__entry__
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_971_to_assign_stmt_977__exit__
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/if_stmt_959_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/if_stmt_959_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_971_to_assign_stmt_977/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_971_to_assign_stmt_977/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_965_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_965_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_965_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_965_PhiAck/$entry
      -- 
    else_choice_transition_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_959_branch_ack_0, ack => convolution3D_CP_1120_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	291 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_update_start_
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Update/cr
      -- 
    ra_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1008_inst_ack_0, ack => convolution3D_CP_1120_elements(131)); -- 
    cr_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(131), ack => RPIPE_maxpool_input_pipe_1008_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Sample/rr
      -- 
    ca_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1008_inst_ack_1, ack => convolution3D_CP_1120_elements(132)); -- 
    rr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(132), ack => type_cast_1012_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Sample/ra
      -- 
    ra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1012_inst_ack_0, ack => convolution3D_CP_1120_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	291 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Update/ca
      -- 
    ca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1012_inst_ack_1, ack => convolution3D_CP_1120_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	291 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Sample/ra
      -- 
    ra_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1027_inst_ack_0, ack => convolution3D_CP_1120_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	291 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Update/ca
      -- 
    ca_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1027_inst_ack_1, ack => convolution3D_CP_1120_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033__exit__
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1034__entry__
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1034_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1034_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1034_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1034_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_436/R_cmpx_xi_1035_place
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1034_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1034_else_link/$entry
      -- 
    branch_req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(137), ack => if_stmt_1034_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(134) & convolution3D_CP_1120_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	281 
    -- CP-element group 138: 	282 
    -- CP-element group 138: 	284 
    -- CP-element group 138: 	285 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_436/if_stmt_1034_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_436/if_stmt_1034_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/$entry
      -- 
    if_choice_transition_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1034_branch_ack_1, ack => convolution3D_CP_1120_elements(138)); -- 
    rr_3429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_986_inst_req_0); -- 
    cr_3434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_986_inst_req_1); -- 
    cr_3457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_993_inst_req_1); -- 
    rr_3452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_993_inst_req_0); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	292 
    -- CP-element group 139: 	293 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Update/cr
      -- CP-element group 139: 	 branch_block_stmt_436/if_stmt_1034_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_436/if_stmt_1034_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- 
    else_choice_transition_2228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1034_branch_ack_0, ack => convolution3D_CP_1120_elements(139)); -- 
    rr_3488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => type_cast_1044_inst_req_0); -- 
    cr_3493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => type_cast_1044_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	295 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_sample_complete
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Sample/ack
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1073_index_offset_ack_0, ack => convolution3D_CP_1120_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	295 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_request/req
      -- 
    ack_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1073_index_offset_ack_1, ack => convolution3D_CP_1120_elements(141)); -- 
    req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(141), ack => addr_of_1074_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_request/$exit
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_request/ack
      -- 
    ack_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1074_final_reg_ack_0, ack => convolution3D_CP_1120_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	295 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/ptr_deref_1077_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/ptr_deref_1077_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/ptr_deref_1077_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/ptr_deref_1077_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/word_access_start/word_0/rr
      -- 
    ack_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1074_final_reg_ack_1, ack => convolution3D_CP_1120_elements(143)); -- 
    rr_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(143), ack => ptr_deref_1077_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Sample/word_access_start/word_0/ra
      -- 
    ra_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1077_store_0_ack_0, ack => convolution3D_CP_1120_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	295 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/word_access_complete/word_0/ca
      -- 
    ca_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1077_store_0_ack_1, ack => convolution3D_CP_1120_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	140 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	296 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079__exit__
      -- CP-element group 146: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/$exit
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(140) & convolution3D_CP_1120_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	296 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Sample/ra
      -- 
    ra_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1084_inst_ack_0, ack => convolution3D_CP_1120_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	296 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	155 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Update/ca
      -- 
    ca_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1084_inst_ack_1, ack => convolution3D_CP_1120_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	296 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Sample/ra
      -- 
    ra_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1088_inst_ack_0, ack => convolution3D_CP_1120_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	296 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	155 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Update/ca
      -- 
    ca_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1088_inst_ack_1, ack => convolution3D_CP_1120_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	296 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Sample/ra
      -- 
    ra_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1092_inst_ack_0, ack => convolution3D_CP_1120_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	296 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Update/ca
      -- 
    ca_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1092_inst_ack_1, ack => convolution3D_CP_1120_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	296 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Sample/ra
      -- 
    ra_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1096_inst_ack_0, ack => convolution3D_CP_1120_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	296 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Update/ca
      -- 
    ca_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1096_inst_ack_1, ack => convolution3D_CP_1120_elements(154)); -- 
    -- CP-element group 155:  branch  join  transition  place  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	148 
    -- CP-element group 155: 	150 
    -- CP-element group 155: 	152 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (10) 
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133__exit__
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1134__entry__
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/$exit
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1134_dead_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1134_eval_test/$entry
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1134_eval_test/$exit
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1134_eval_test/branch_req
      -- CP-element group 155: 	 branch_block_stmt_436/R_cmp161317_1135_place
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1134_if_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1134_else_link/$entry
      -- 
    branch_req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(155), ack => if_stmt_1134_branch_req_0); -- 
    convolution3D_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(148) & convolution3D_CP_1120_elements(150) & convolution3D_CP_1120_elements(152) & convolution3D_CP_1120_elements(154);
      gj_convolution3D_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: 	159 
    -- CP-element group 156: 	160 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	162 
    -- CP-element group 156: 	163 
    -- CP-element group 156: 	164 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	168 
    -- CP-element group 156: 	170 
    -- CP-element group 156:  members (42) 
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1140__exit__
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211__entry__
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1140_PhiReqMerge
      -- CP-element group 156: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1140_PhiAck/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1140_PhiAck/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1140_PhiAck/dummy
      -- CP-element group 156: 	 branch_block_stmt_436/if_stmt_1134_if_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/if_stmt_1134_if_link/if_choice_transition
      -- CP-element group 156: 	 branch_block_stmt_436/ifx_xend_bbx_xnph
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Update/cr
      -- 
    if_choice_transition_2401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1134_branch_ack_1, ack => convolution3D_CP_1120_elements(156)); -- 
    rr_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1155_inst_req_0); -- 
    cr_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1155_inst_req_1); -- 
    rr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1159_inst_req_0); -- 
    cr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1159_inst_req_1); -- 
    rr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1168_inst_req_0); -- 
    cr_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1168_inst_req_1); -- 
    rr_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1177_inst_req_0); -- 
    cr_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1177_inst_req_1); -- 
    cr_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1186_inst_req_1); -- 
    cr_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1191_inst_req_1); -- 
    -- CP-element group 157:  transition  place  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	306 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_436/if_stmt_1134_else_link/$exit
      -- CP-element group 157: 	 branch_block_stmt_436/if_stmt_1134_else_link/else_choice_transition
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$entry
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1408/$entry
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/$entry
      -- 
    else_choice_transition_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1134_branch_ack_0, ack => convolution3D_CP_1120_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Sample/ra
      -- 
    ra_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1155_inst_ack_0, ack => convolution3D_CP_1120_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	156 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	166 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1155_Update/ca
      -- 
    ca_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1155_inst_ack_1, ack => convolution3D_CP_1120_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	156 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Sample/ra
      -- 
    ra_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_0, ack => convolution3D_CP_1120_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	166 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1159_Update/ca
      -- 
    ca_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_1, ack => convolution3D_CP_1120_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	156 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Sample/ra
      -- 
    ra_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_0, ack => convolution3D_CP_1120_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	156 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1168_Update/ca
      -- 
    ca_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_1, ack => convolution3D_CP_1120_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Sample/ra
      -- 
    ra_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_0, ack => convolution3D_CP_1120_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1177_Update/ca
      -- 
    ca_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_1, ack => convolution3D_CP_1120_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	159 
    -- CP-element group 166: 	161 
    -- CP-element group 166: 	163 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Sample/rr
      -- 
    rr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(166), ack => type_cast_1186_inst_req_0); -- 
    convolution3D_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(159) & convolution3D_CP_1120_elements(161) & convolution3D_CP_1120_elements(163) & convolution3D_CP_1120_elements(165);
      gj_convolution3D_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Sample/ra
      -- 
    ra_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_0, ack => convolution3D_CP_1120_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	156 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1186_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Sample/rr
      -- 
    ca_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_1, ack => convolution3D_CP_1120_elements(168)); -- 
    rr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(168), ack => type_cast_1191_inst_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Sample/ra
      -- 
    ra_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_0, ack => convolution3D_CP_1120_elements(169)); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	156 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	297 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211__exit__
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1214/$entry
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/$entry
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/$exit
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1146_to_assign_stmt_1211/type_cast_1191_Update/ca
      -- 
    ca_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_1, ack => convolution3D_CP_1120_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	302 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	210 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_sample_complete
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Sample/ack
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Sample/$exit
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1226_index_offset_ack_0, ack => convolution3D_CP_1120_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	302 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (11) 
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_request/$entry
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_request/req
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_offset_calculated
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1226_index_offset_ack_1, ack => convolution3D_CP_1120_elements(172)); -- 
    req_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(172), ack => addr_of_1227_final_reg_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_request/$exit
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_request/ack
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_sample_completed_
      -- 
    ack_2538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1227_final_reg_ack_0, ack => convolution3D_CP_1120_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	302 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	207 
    -- CP-element group 174:  members (19) 
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_complete/ack
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_word_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_address_resized
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_addr_resize/$entry
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_addr_resize/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_addr_resize/base_resize_req
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_addr_resize/base_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_base_plus_offset/sum_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_word_addrgen/$entry
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_word_addrgen/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_word_addrgen/root_register_req
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_word_addrgen/root_register_ack
      -- 
    ack_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1227_final_reg_ack_1, ack => convolution3D_CP_1120_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	302 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_update_start_
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_sample_completed_
      -- 
    ra_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1230_inst_ack_0, ack => convolution3D_CP_1120_elements(175)); -- 
    cr_2556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(175), ack => RPIPE_maxpool_input_pipe_1230_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_update_completed_
      -- 
    ca_2557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1230_inst_ack_1, ack => convolution3D_CP_1120_elements(176)); -- 
    rr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(176), ack => type_cast_1234_inst_req_0); -- 
    rr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(176), ack => RPIPE_maxpool_input_pipe_1243_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Sample/$exit
      -- 
    ra_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_0, ack => convolution3D_CP_1120_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	302 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	207 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Update/ca
      -- 
    ca_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_1, ack => convolution3D_CP_1120_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_update_start_
      -- 
    ra_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1243_inst_ack_0, ack => convolution3D_CP_1120_elements(179)); -- 
    cr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(179), ack => RPIPE_maxpool_input_pipe_1243_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1243_Update/ca
      -- 
    ca_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1243_inst_ack_1, ack => convolution3D_CP_1120_elements(180)); -- 
    rr_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => type_cast_1247_inst_req_0); -- 
    rr_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => RPIPE_maxpool_input_pipe_1261_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_sample_completed_
      -- 
    ra_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_0, ack => convolution3D_CP_1120_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	302 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	207 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_update_completed_
      -- 
    ca_2599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_1, ack => convolution3D_CP_1120_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_update_start_
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_sample_completed_
      -- 
    ra_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1261_inst_ack_0, ack => convolution3D_CP_1120_elements(183)); -- 
    cr_2612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(183), ack => RPIPE_maxpool_input_pipe_1261_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1261_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Sample/rr
      -- 
    ca_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1261_inst_ack_1, ack => convolution3D_CP_1120_elements(184)); -- 
    rr_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(184), ack => type_cast_1265_inst_req_0); -- 
    rr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(184), ack => RPIPE_maxpool_input_pipe_1279_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Sample/$exit
      -- 
    ra_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_0, ack => convolution3D_CP_1120_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	302 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	207 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Update/ca
      -- 
    ca_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_1, ack => convolution3D_CP_1120_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_update_start_
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Sample/$exit
      -- 
    ra_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1279_inst_ack_0, ack => convolution3D_CP_1120_elements(187)); -- 
    cr_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => RPIPE_maxpool_input_pipe_1279_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1279_Update/$exit
      -- 
    ca_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1279_inst_ack_1, ack => convolution3D_CP_1120_elements(188)); -- 
    rr_2649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(188), ack => type_cast_1283_inst_req_0); -- 
    rr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(188), ack => RPIPE_maxpool_input_pipe_1297_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_sample_completed_
      -- 
    ra_2650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_0, ack => convolution3D_CP_1120_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	302 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	207 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_update_completed_
      -- 
    ca_2655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_1, ack => convolution3D_CP_1120_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_update_start_
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Sample/ra
      -- 
    ra_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1297_inst_ack_0, ack => convolution3D_CP_1120_elements(191)); -- 
    cr_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(191), ack => RPIPE_maxpool_input_pipe_1297_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1297_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_sample_start_
      -- 
    ca_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1297_inst_ack_1, ack => convolution3D_CP_1120_elements(192)); -- 
    rr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(192), ack => type_cast_1301_inst_req_0); -- 
    rr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(192), ack => RPIPE_maxpool_input_pipe_1315_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_sample_completed_
      -- 
    ra_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_0, ack => convolution3D_CP_1120_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	302 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	207 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Update/$exit
      -- 
    ca_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_1, ack => convolution3D_CP_1120_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Update/cr
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_update_start_
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_sample_completed_
      -- 
    ra_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1315_inst_ack_0, ack => convolution3D_CP_1120_elements(195)); -- 
    cr_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(195), ack => RPIPE_maxpool_input_pipe_1315_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1315_update_completed_
      -- 
    ca_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1315_inst_ack_1, ack => convolution3D_CP_1120_elements(196)); -- 
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(196), ack => type_cast_1319_inst_req_0); -- 
    rr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(196), ack => RPIPE_maxpool_input_pipe_1333_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Sample/ra
      -- 
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1319_inst_ack_0, ack => convolution3D_CP_1120_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	302 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	207 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Update/$exit
      -- 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1319_inst_ack_1, ack => convolution3D_CP_1120_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_update_start_
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Update/cr
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Sample/ra
      -- 
    ra_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1333_inst_ack_0, ack => convolution3D_CP_1120_elements(199)); -- 
    cr_2724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(199), ack => RPIPE_maxpool_input_pipe_1333_inst_req_1); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1333_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Sample/rr
      -- 
    ca_2725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1333_inst_ack_1, ack => convolution3D_CP_1120_elements(200)); -- 
    rr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(200), ack => type_cast_1337_inst_req_0); -- 
    rr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(200), ack => RPIPE_maxpool_input_pipe_1351_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Sample/ra
      -- 
    ra_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1337_inst_ack_0, ack => convolution3D_CP_1120_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	302 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Update/ca
      -- 
    ca_2739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1337_inst_ack_1, ack => convolution3D_CP_1120_elements(202)); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_update_start_
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Update/cr
      -- 
    ra_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1351_inst_ack_0, ack => convolution3D_CP_1120_elements(203)); -- 
    cr_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(203), ack => RPIPE_maxpool_input_pipe_1351_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1351_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Sample/rr
      -- 
    ca_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1351_inst_ack_1, ack => convolution3D_CP_1120_elements(204)); -- 
    rr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(204), ack => type_cast_1355_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Sample/ra
      -- 
    ra_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1355_inst_ack_0, ack => convolution3D_CP_1120_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	302 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Update/ca
      -- 
    ca_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1355_inst_ack_1, ack => convolution3D_CP_1120_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	174 
    -- CP-element group 207: 	178 
    -- CP-element group 207: 	182 
    -- CP-element group 207: 	186 
    -- CP-element group 207: 	190 
    -- CP-element group 207: 	194 
    -- CP-element group 207: 	198 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/ptr_deref_1363_Split/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/ptr_deref_1363_Split/$exit
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/ptr_deref_1363_Split/split_req
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/ptr_deref_1363_Split/split_ack
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/word_access_start/word_0/rr
      -- 
    rr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(207), ack => ptr_deref_1363_store_0_req_0); -- 
    convolution3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(174) & convolution3D_CP_1120_elements(178) & convolution3D_CP_1120_elements(182) & convolution3D_CP_1120_elements(186) & convolution3D_CP_1120_elements(190) & convolution3D_CP_1120_elements(194) & convolution3D_CP_1120_elements(198) & convolution3D_CP_1120_elements(202) & convolution3D_CP_1120_elements(206);
      gj_convolution3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/word_access_start/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/word_access_start/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Sample/word_access_start/word_0/ra
      -- 
    ra_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1363_store_0_ack_0, ack => convolution3D_CP_1120_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	302 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/word_access_complete/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/word_access_complete/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/word_access_complete/word_0/ca
      -- 
    ca_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1363_store_0_ack_1, ack => convolution3D_CP_1120_elements(209)); -- 
    -- CP-element group 210:  branch  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	171 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (10) 
      -- CP-element group 210: 	 branch_block_stmt_436/R_exitcond_1378_place
      -- CP-element group 210: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376__exit__
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1377__entry__
      -- CP-element group 210: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/$exit
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1377_dead_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1377_eval_test/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1377_eval_test/$exit
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1377_eval_test/branch_req
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1377_if_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1377_else_link/$entry
      -- 
    branch_req_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(210), ack => if_stmt_1377_branch_req_0); -- 
    convolution3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(171) & convolution3D_CP_1120_elements(209);
      gj_convolution3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	303 
    -- CP-element group 211: 	304 
    -- CP-element group 211:  members (24) 
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1383_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1383__exit__
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1390_to_assign_stmt_1405__entry__
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1390_to_assign_stmt_1405__exit__
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 211: 	 branch_block_stmt_436/if_stmt_1377_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/if_stmt_1377_if_link/if_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1390_to_assign_stmt_1405/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1390_to_assign_stmt_1405/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Update/cr
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1383_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1383_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1383_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- 
    if_choice_transition_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1377_branch_ack_1, ack => convolution3D_CP_1120_elements(211)); -- 
    cr_3601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => type_cast_1411_inst_req_1); -- 
    rr_3596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => type_cast_1411_inst_req_0); -- 
    -- CP-element group 212:  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	298 
    -- CP-element group 212: 	299 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/if_stmt_1377_else_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_436/if_stmt_1377_else_link/else_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1377_branch_ack_0, ack => convolution3D_CP_1120_elements(212)); -- 
    rr_3553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_1220_inst_req_0); -- 
    cr_3558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_1220_inst_req_1); -- 
    -- CP-element group 213:  transition  place  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	308 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	327 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_436/forx_xend215_ifx_xend227
      -- CP-element group 213: 	 branch_block_stmt_436/if_stmt_1428_if_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_436/if_stmt_1428_if_link/if_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_436/forx_xend215_ifx_xend227_PhiReq/$exit
      -- CP-element group 213: 	 branch_block_stmt_436/forx_xend215_ifx_xend227_PhiReq/$entry
      -- 
    if_choice_transition_2855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1428_branch_ack_1, ack => convolution3D_CP_1120_elements(213)); -- 
    -- CP-element group 214:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	308 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (18) 
      -- CP-element group 214: 	 branch_block_stmt_436/forx_xend215_bbx_xnphx_xi294
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1434_PhiReqMerge
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1434__exit__
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450__entry__
      -- CP-element group 214: 	 branch_block_stmt_436/forx_xend215_bbx_xnphx_xi294_PhiReq/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/forx_xend215_bbx_xnphx_xi294_PhiReq/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1434_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1434_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1434_PhiAck/dummy
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1428_else_link/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1428_else_link/else_choice_transition
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_update_start_
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Update/cr
      -- 
    else_choice_transition_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1428_branch_ack_0, ack => convolution3D_CP_1120_elements(214)); -- 
    rr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(214), ack => type_cast_1443_inst_req_0); -- 
    cr_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(214), ack => type_cast_1443_inst_req_1); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Sample/ra
      -- 
    ra_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1443_inst_ack_0, ack => convolution3D_CP_1120_elements(215)); -- 
    -- CP-element group 216:  fork  transition  place  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	309 
    -- CP-element group 216: 	310 
    -- CP-element group 216:  members (11) 
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450__exit__
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1440_to_assign_stmt_1450/type_cast_1443_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/$entry
      -- 
    ca_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1443_inst_ack_1, ack => convolution3D_CP_1120_elements(216)); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	322 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_update_start_
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Update/cr
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1481_inst_ack_0, ack => convolution3D_CP_1120_elements(217)); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(217), ack => RPIPE_maxpool_input_pipe_1481_inst_req_1); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Sample/rr
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1481_inst_ack_1, ack => convolution3D_CP_1120_elements(218)); -- 
    rr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => type_cast_1485_inst_req_0); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Sample/ra
      -- 
    ra_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1485_inst_ack_0, ack => convolution3D_CP_1120_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	322 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Update/ca
      -- 
    ca_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1485_inst_ack_1, ack => convolution3D_CP_1120_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	322 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Sample/ra
      -- 
    ra_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1500_inst_ack_0, ack => convolution3D_CP_1120_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	322 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Update/ca
      -- 
    ca_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1500_inst_ack_1, ack => convolution3D_CP_1120_elements(222)); -- 
    -- CP-element group 223:  branch  join  transition  place  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (10) 
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506__exit__
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1507__entry__
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/$exit
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1507_dead_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1507_eval_test/$entry
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1507_eval_test/$exit
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1507_eval_test/branch_req
      -- CP-element group 223: 	 branch_block_stmt_436/R_cmpx_xi302_1508_place
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1507_if_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1507_else_link/$entry
      -- 
    branch_req_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(223), ack => if_stmt_1507_branch_req_0); -- 
    convolution3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(220) & convolution3D_CP_1120_elements(222);
      gj_convolution3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	312 
    -- CP-element group 224: 	313 
    -- CP-element group 224: 	315 
    -- CP-element group 224: 	316 
    -- CP-element group 224:  members (20) 
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/if_stmt_1507_if_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_436/if_stmt_1507_if_link/if_choice_transition
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1507_branch_ack_1, ack => convolution3D_CP_1120_elements(224)); -- 
    rr_3669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1459_inst_req_0); -- 
    cr_3674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1459_inst_req_1); -- 
    rr_3692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1466_inst_req_0); -- 
    cr_3697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1466_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  place  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	323 
    -- CP-element group 225: 	324 
    -- CP-element group 225:  members (12) 
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/if_stmt_1507_else_link/$exit
      -- CP-element group 225: 	 branch_block_stmt_436/if_stmt_1507_else_link/else_choice_transition
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1507_branch_ack_0, ack => convolution3D_CP_1120_elements(225)); -- 
    rr_3728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(225), ack => type_cast_1517_inst_req_0); -- 
    cr_3733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(225), ack => type_cast_1517_inst_req_1); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	326 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	232 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_sample_complete
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Sample/ack
      -- 
    ack_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1546_index_offset_ack_0, ack => convolution3D_CP_1120_elements(226)); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	326 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (11) 
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_offset_calculated
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Update/ack
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_base_plus_offset/$entry
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_base_plus_offset/$exit
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_base_plus_offset/sum_rename_req
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_base_plus_offset/sum_rename_ack
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_request/$entry
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_request/req
      -- 
    ack_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1546_index_offset_ack_1, ack => convolution3D_CP_1120_elements(227)); -- 
    req_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(227), ack => addr_of_1547_final_reg_req_0); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_request/$exit
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_request/ack
      -- 
    ack_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1547_final_reg_ack_0, ack => convolution3D_CP_1120_elements(228)); -- 
    -- CP-element group 229:  join  fork  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	326 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (28) 
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_complete/ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_word_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_root_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_address_resized
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_addr_resize/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_addr_resize/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_addr_resize/base_resize_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_addr_resize/base_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_plus_offset/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_plus_offset/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_plus_offset/sum_rename_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_base_plus_offset/sum_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_word_addrgen/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_word_addrgen/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_word_addrgen/root_register_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_word_addrgen/root_register_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/ptr_deref_1550_Split/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/ptr_deref_1550_Split/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/ptr_deref_1550_Split/split_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/ptr_deref_1550_Split/split_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/word_access_start/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/word_access_start/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/word_access_start/word_0/rr
      -- 
    ack_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1547_final_reg_ack_1, ack => convolution3D_CP_1120_elements(229)); -- 
    rr_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(229), ack => ptr_deref_1550_store_0_req_0); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Sample/word_access_start/word_0/ra
      -- 
    ra_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1550_store_0_ack_0, ack => convolution3D_CP_1120_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	326 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (5) 
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/word_access_complete/word_0/ca
      -- 
    ca_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1550_store_0_ack_1, ack => convolution3D_CP_1120_elements(231)); -- 
    -- CP-element group 232:  join  transition  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	226 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	327 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552__exit__
      -- CP-element group 232: 	 branch_block_stmt_436/getRemainingElementsx_xexit311_ifx_xend227
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/$exit
      -- CP-element group 232: 	 branch_block_stmt_436/getRemainingElementsx_xexit311_ifx_xend227_PhiReq/$exit
      -- CP-element group 232: 	 branch_block_stmt_436/getRemainingElementsx_xexit311_ifx_xend227_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(226) & convolution3D_CP_1120_elements(231);
      gj_convolution3D_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	327 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Sample/cra
      -- 
    cra_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1557_call_ack_0, ack => convolution3D_CP_1120_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	327 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	237 
    -- CP-element group 234: 	239 
    -- CP-element group 234: 	240 
    -- CP-element group 234: 	241 
    -- CP-element group 234: 	242 
    -- CP-element group 234: 	243 
    -- CP-element group 234: 	244 
    -- CP-element group 234:  members (31) 
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1557__exit__
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621__entry__
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1557/$exit
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Update/cca
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_update_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_update_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_update_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Update/cr
      -- 
    cca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1557_call_ack_1, ack => convolution3D_CP_1120_elements(234)); -- 
    req_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => WPIPE_num_out_pipe_1569_inst_req_0); -- 
    req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => WPIPE_maxpool_output_pipe_1572_inst_req_0); -- 
    rr_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1596_inst_req_0); -- 
    cr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1596_inst_req_1); -- 
    rr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1606_inst_req_0); -- 
    cr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1606_inst_req_1); -- 
    rr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1615_inst_req_0); -- 
    cr_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1615_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_update_start_
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Update/req
      -- 
    ack_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1569_inst_ack_0, ack => convolution3D_CP_1120_elements(235)); -- 
    req_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(235), ack => WPIPE_num_out_pipe_1569_inst_req_1); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	245 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_num_out_pipe_1569_Update/ack
      -- 
    ack_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1569_inst_ack_1, ack => convolution3D_CP_1120_elements(236)); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	234 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_update_start_
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Update/req
      -- 
    ack_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1572_inst_ack_0, ack => convolution3D_CP_1120_elements(237)); -- 
    req_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(237), ack => WPIPE_maxpool_output_pipe_1572_inst_req_1); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	245 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/WPIPE_maxpool_output_pipe_1572_Update/ack
      -- 
    ack_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1572_inst_ack_1, ack => convolution3D_CP_1120_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	234 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Sample/ra
      -- 
    ra_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1596_inst_ack_0, ack => convolution3D_CP_1120_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	234 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	245 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1596_Update/ca
      -- 
    ca_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1596_inst_ack_1, ack => convolution3D_CP_1120_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	234 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Sample/ra
      -- 
    ra_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_0, ack => convolution3D_CP_1120_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	234 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	245 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1606_Update/ca
      -- 
    ca_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_1, ack => convolution3D_CP_1120_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	234 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Sample/ra
      -- 
    ra_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_0, ack => convolution3D_CP_1120_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	234 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/type_cast_1615_Update/ca
      -- 
    ca_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_1, ack => convolution3D_CP_1120_elements(244)); -- 
    -- CP-element group 245:  join  transition  place  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	236 
    -- CP-element group 245: 	238 
    -- CP-element group 245: 	240 
    -- CP-element group 245: 	242 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	328 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621__exit__
      -- CP-element group 245: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody
      -- CP-element group 245: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$entry
      -- CP-element group 245: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1624/$entry
      -- CP-element group 245: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1563_to_assign_stmt_1621/$exit
      -- 
    convolution3D_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(236) & convolution3D_CP_1120_elements(238) & convolution3D_CP_1120_elements(240) & convolution3D_CP_1120_elements(242) & convolution3D_CP_1120_elements(244);
      gj_convolution3D_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	333 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Sample/ra
      -- 
    ra_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_0, ack => convolution3D_CP_1120_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	333 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	250 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Update/ca
      -- 
    ca_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_1, ack => convolution3D_CP_1120_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	333 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Sample/ra
      -- 
    ra_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1648_inst_ack_0, ack => convolution3D_CP_1120_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	333 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Update/ca
      -- 
    ca_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1648_inst_ack_1, ack => convolution3D_CP_1120_elements(249)); -- 
    -- CP-element group 250:  join  transition  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	247 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Sample/crr
      -- 
    crr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(250), ack => call_stmt_1652_call_req_0); -- 
    convolution3D_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(247) & convolution3D_CP_1120_elements(249);
      gj_convolution3D_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Sample/cra
      -- 
    cra_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1652_call_ack_0, ack => convolution3D_CP_1120_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	333 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	255 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Update/cca
      -- 
    cca_3176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1652_call_ack_1, ack => convolution3D_CP_1120_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	333 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Sample/cra
      -- 
    cra_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1659_call_ack_0, ack => convolution3D_CP_1120_elements(253)); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	333 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Update/cca
      -- 
    cca_3190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1659_call_ack_1, ack => convolution3D_CP_1120_elements(254)); -- 
    -- CP-element group 255:  branch  join  transition  place  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	252 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (10) 
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670__exit__
      -- CP-element group 255: 	 branch_block_stmt_436/if_stmt_1671__entry__
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/$exit
      -- CP-element group 255: 	 branch_block_stmt_436/if_stmt_1671_dead_link/$entry
      -- CP-element group 255: 	 branch_block_stmt_436/if_stmt_1671_eval_test/$entry
      -- CP-element group 255: 	 branch_block_stmt_436/if_stmt_1671_eval_test/$exit
      -- CP-element group 255: 	 branch_block_stmt_436/if_stmt_1671_eval_test/branch_req
      -- CP-element group 255: 	 branch_block_stmt_436/R_exitcond5_1672_place
      -- CP-element group 255: 	 branch_block_stmt_436/if_stmt_1671_if_link/$entry
      -- CP-element group 255: 	 branch_block_stmt_436/if_stmt_1671_else_link/$entry
      -- 
    branch_req_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(255), ack => if_stmt_1671_branch_req_0); -- 
    convolution3D_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(252) & convolution3D_CP_1120_elements(254);
      gj_convolution3D_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: 	259 
    -- CP-element group 256:  members (18) 
      -- CP-element group 256: 	 branch_block_stmt_436/merge_stmt_1677__exit__
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682__entry__
      -- CP-element group 256: 	 branch_block_stmt_436/merge_stmt_1677_PhiReqMerge
      -- CP-element group 256: 	 branch_block_stmt_436/if_stmt_1671_if_link/$exit
      -- CP-element group 256: 	 branch_block_stmt_436/if_stmt_1671_if_link/if_choice_transition
      -- CP-element group 256: 	 branch_block_stmt_436/whilex_xbody_whilex_xend
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682/$entry
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_update_start_
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Sample/rr
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Update/cr
      -- CP-element group 256: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 256: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 256: 	 branch_block_stmt_436/merge_stmt_1677_PhiAck/$entry
      -- CP-element group 256: 	 branch_block_stmt_436/merge_stmt_1677_PhiAck/$exit
      -- CP-element group 256: 	 branch_block_stmt_436/merge_stmt_1677_PhiAck/dummy
      -- 
    if_choice_transition_3203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1671_branch_ack_1, ack => convolution3D_CP_1120_elements(256)); -- 
    rr_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(256), ack => type_cast_1681_inst_req_0); -- 
    cr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(256), ack => type_cast_1681_inst_req_1); -- 
    -- CP-element group 257:  fork  transition  place  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	329 
    -- CP-element group 257: 	330 
    -- CP-element group 257:  members (12) 
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/cr
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/rr
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1671_else_link/$exit
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1671_else_link/else_choice_transition
      -- CP-element group 257: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody
      -- 
    else_choice_transition_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1671_branch_ack_0, ack => convolution3D_CP_1120_elements(257)); -- 
    cr_3786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(257), ack => type_cast_1627_inst_req_1); -- 
    rr_3781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(257), ack => type_cast_1627_inst_req_0); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Sample/ra
      -- 
    ra_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1681_inst_ack_0, ack => convolution3D_CP_1120_elements(258)); -- 
    -- CP-element group 259:  fork  transition  place  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	256 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259: 	261 
    -- CP-element group 259: 	263 
    -- CP-element group 259:  members (16) 
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1682__exit__
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698__entry__
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1682/$exit
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1682/type_cast_1681_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_update_start_
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Sample/crr
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Update/ccr
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_update_start_
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Update/cr
      -- 
    ca_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1681_inst_ack_1, ack => convolution3D_CP_1120_elements(259)); -- 
    crr_3237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(259), ack => call_stmt_1685_call_req_0); -- 
    ccr_3242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(259), ack => call_stmt_1685_call_req_1); -- 
    cr_3256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(259), ack => type_cast_1689_inst_req_1); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Sample/cra
      -- 
    cra_3238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1685_call_ack_0, ack => convolution3D_CP_1120_elements(260)); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/call_stmt_1685_Update/cca
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Sample/rr
      -- 
    cca_3243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1685_call_ack_1, ack => convolution3D_CP_1120_elements(261)); -- 
    rr_3251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(261), ack => type_cast_1689_inst_req_0); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Sample/ra
      -- 
    ra_3252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1689_inst_ack_0, ack => convolution3D_CP_1120_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	259 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/type_cast_1689_Update/ca
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Sample/req
      -- 
    ca_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1689_inst_ack_1, ack => convolution3D_CP_1120_elements(263)); -- 
    req_3265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(263), ack => WPIPE_elapsed_time_pipe_1696_inst_req_0); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_update_start_
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Sample/ack
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Update/req
      -- 
    ack_3266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1696_inst_ack_0, ack => convolution3D_CP_1120_elements(264)); -- 
    req_3270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(264), ack => WPIPE_elapsed_time_pipe_1696_inst_req_1); -- 
    -- CP-element group 265:  transition  place  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (16) 
      -- CP-element group 265: 	 $exit
      -- CP-element group 265: 	 branch_block_stmt_436/$exit
      -- CP-element group 265: 	 branch_block_stmt_436/branch_block_stmt_436__exit__
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698__exit__
      -- CP-element group 265: 	 branch_block_stmt_436/return__
      -- CP-element group 265: 	 branch_block_stmt_436/merge_stmt_1701__exit__
      -- CP-element group 265: 	 branch_block_stmt_436/merge_stmt_1701_PhiReqMerge
      -- CP-element group 265: 	 branch_block_stmt_436/merge_stmt_1701_PhiAck/$entry
      -- CP-element group 265: 	 branch_block_stmt_436/merge_stmt_1701_PhiAck/$exit
      -- CP-element group 265: 	 branch_block_stmt_436/merge_stmt_1701_PhiAck/dummy
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/$exit
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1685_to_assign_stmt_1698/WPIPE_elapsed_time_pipe_1696_Update/ack
      -- CP-element group 265: 	 branch_block_stmt_436/return___PhiReq/$entry
      -- CP-element group 265: 	 branch_block_stmt_436/return___PhiReq/$exit
      -- 
    ack_3271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1696_inst_ack_1, ack => convolution3D_CP_1120_elements(265)); -- 
    -- CP-element group 266:  transition  output  delay-element  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	86 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	270 
    -- CP-element group 266:  members (5) 
      -- CP-element group 266: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/$exit
      -- CP-element group 266: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_745/$exit
      -- CP-element group 266: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/$exit
      -- CP-element group 266: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_749_konst_delay_trans
      -- CP-element group 266: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_req
      -- 
    phi_stmt_745_req_3294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_745_req_3294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(266), ack => phi_stmt_745_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(266) is a control-delay.
    cp_element_266_delay: control_delay_element  generic map(name => " 266_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(86), ack => convolution3D_CP_1120_elements(266), clk => clk, reset =>reset);
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	128 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (2) 
      -- CP-element group 267: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Sample/ra
      -- 
    ra_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => convolution3D_CP_1120_elements(267)); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	128 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (2) 
      -- CP-element group 268: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/Update/ca
      -- 
    ca_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_1, ack => convolution3D_CP_1120_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/$exit
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/$exit
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/$exit
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_sources/type_cast_751/SplitProtocol/$exit
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_745/phi_stmt_745_req
      -- 
    phi_stmt_745_req_3320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_745_req_3320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(269), ack => phi_stmt_745_req_1); -- 
    convolution3D_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(267) & convolution3D_CP_1120_elements(268);
      gj_convolution3D_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  merge  transition  place  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	266 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_436/merge_stmt_744_PhiReqMerge
      -- CP-element group 270: 	 branch_block_stmt_436/merge_stmt_744_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(270) <= OrReduce(convolution3D_CP_1120_elements(266) & convolution3D_CP_1120_elements(269));
    -- CP-element group 271:  fork  transition  place  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	87 
    -- CP-element group 271: 	88 
    -- CP-element group 271: 	90 
    -- CP-element group 271: 	91 
    -- CP-element group 271: 	94 
    -- CP-element group 271: 	98 
    -- CP-element group 271: 	102 
    -- CP-element group 271: 	106 
    -- CP-element group 271: 	110 
    -- CP-element group 271: 	114 
    -- CP-element group 271: 	118 
    -- CP-element group 271: 	122 
    -- CP-element group 271: 	125 
    -- CP-element group 271:  members (56) 
      -- CP-element group 271: 	 branch_block_stmt_436/merge_stmt_744__exit__
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907__entry__
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_resized_1
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_scaled_1
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_computed_1
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_resize_1/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_resize_1/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_resize_1/index_resize_req
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_resize_1/index_resize_ack
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_scale_1/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_scale_1/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_scale_1/scale_rename_req
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_index_scale_1/scale_rename_ack
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_update_start
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Sample/req
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/array_obj_ref_757_final_index_sum_regn_Update/req
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_complete/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/addr_of_758_complete/req
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/RPIPE_maxpool_input_pipe_761_Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_765_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_778_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_796_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_814_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_832_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_850_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_868_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/type_cast_886_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_update_start_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/word_access_complete/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/word_access_complete/word_0/$entry
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_759_to_assign_stmt_907/ptr_deref_894_Update/word_access_complete/word_0/cr
      -- CP-element group 271: 	 branch_block_stmt_436/merge_stmt_744_PhiAck/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/merge_stmt_744_PhiAck/phi_stmt_745_ack
      -- 
    phi_stmt_745_ack_3325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_745_ack_0, ack => convolution3D_CP_1120_elements(271)); -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => array_obj_ref_757_index_offset_req_0); -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => array_obj_ref_757_index_offset_req_1); -- 
    req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => addr_of_758_final_reg_req_1); -- 
    rr_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => RPIPE_maxpool_input_pipe_761_inst_req_0); -- 
    cr_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_765_inst_req_1); -- 
    cr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_778_inst_req_1); -- 
    cr_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_796_inst_req_1); -- 
    cr_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_814_inst_req_1); -- 
    cr_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_832_inst_req_1); -- 
    cr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_850_inst_req_1); -- 
    cr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_868_inst_req_1); -- 
    cr_2068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => type_cast_886_inst_req_1); -- 
    cr_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => ptr_deref_894_store_0_req_1); -- 
    -- CP-element group 272:  transition  output  delay-element  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	76 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	276 
    -- CP-element group 272:  members (5) 
      -- CP-element group 272: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/$exit
      -- CP-element group 272: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_939/$exit
      -- CP-element group 272: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_945_konst_delay_trans
      -- CP-element group 272: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_req
      -- CP-element group 272: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_939_req_3348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_939_req_3348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(272), ack => phi_stmt_939_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(272) is a control-delay.
    cp_element_272_delay: control_delay_element  generic map(name => " 272_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(76), ack => convolution3D_CP_1120_elements(272), clk => clk, reset =>reset);
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	127 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Sample/ra
      -- 
    ra_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_942_inst_ack_0, ack => convolution3D_CP_1120_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	127 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Update/ca
      -- CP-element group 274: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/Update/$exit
      -- 
    ca_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_942_inst_ack_1, ack => convolution3D_CP_1120_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_req
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/$exit
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/$exit
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/$exit
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_939/phi_stmt_939_sources/type_cast_942/SplitProtocol/$exit
      -- 
    phi_stmt_939_req_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_939_req_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(275), ack => phi_stmt_939_req_0); -- 
    convolution3D_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(273) & convolution3D_CP_1120_elements(274);
      gj_convolution3D_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  merge  transition  place  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	272 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (2) 
      -- CP-element group 276: 	 branch_block_stmt_436/merge_stmt_938_PhiAck/$entry
      -- CP-element group 276: 	 branch_block_stmt_436/merge_stmt_938_PhiReqMerge
      -- 
    convolution3D_CP_1120_elements(276) <= OrReduce(convolution3D_CP_1120_elements(272) & convolution3D_CP_1120_elements(275));
    -- CP-element group 277:  branch  transition  place  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	129 
    -- CP-element group 277: 	130 
    -- CP-element group 277:  members (15) 
      -- CP-element group 277: 	 branch_block_stmt_436/merge_stmt_938__exit__
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_952_to_assign_stmt_958__entry__
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_952_to_assign_stmt_958__exit__
      -- CP-element group 277: 	 branch_block_stmt_436/if_stmt_959__entry__
      -- CP-element group 277: 	 branch_block_stmt_436/merge_stmt_938_PhiAck/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/merge_stmt_938_PhiAck/phi_stmt_939_ack
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_952_to_assign_stmt_958/$entry
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_952_to_assign_stmt_958/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/if_stmt_959_dead_link/$entry
      -- CP-element group 277: 	 branch_block_stmt_436/if_stmt_959_eval_test/$entry
      -- CP-element group 277: 	 branch_block_stmt_436/if_stmt_959_eval_test/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/if_stmt_959_eval_test/branch_req
      -- CP-element group 277: 	 branch_block_stmt_436/R_tobool_960_place
      -- CP-element group 277: 	 branch_block_stmt_436/if_stmt_959_if_link/$entry
      -- CP-element group 277: 	 branch_block_stmt_436/if_stmt_959_else_link/$entry
      -- 
    phi_stmt_939_ack_3379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_939_ack_0, ack => convolution3D_CP_1120_elements(277)); -- 
    branch_req_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(277), ack => if_stmt_959_branch_req_0); -- 
    -- CP-element group 278:  transition  output  delay-element  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	130 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (4) 
      -- CP-element group 278: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_req
      -- CP-element group 278: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_984_konst_delay_trans
      -- CP-element group 278: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/$exit
      -- CP-element group 278: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/$exit
      -- 
    phi_stmt_980_req_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_980_req_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(278), ack => phi_stmt_980_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(278) is a control-delay.
    cp_element_278_delay: control_delay_element  generic map(name => " 278_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(130), ack => convolution3D_CP_1120_elements(278), clk => clk, reset =>reset);
    -- CP-element group 279:  transition  output  delay-element  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	130 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (4) 
      -- CP-element group 279: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/$exit
      -- CP-element group 279: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_991_konst_delay_trans
      -- CP-element group 279: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_req
      -- 
    phi_stmt_987_req_3410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_987_req_3410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(279), ack => phi_stmt_987_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(279) is a control-delay.
    cp_element_279_delay: control_delay_element  generic map(name => " 279_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(130), ack => convolution3D_CP_1120_elements(279), clk => clk, reset =>reset);
    -- CP-element group 280:  join  transition  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	288 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(278) & convolution3D_CP_1120_elements(279);
      gj_convolution3D_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	138 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Sample/ra
      -- 
    ra_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_986_inst_ack_0, ack => convolution3D_CP_1120_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	138 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (2) 
      -- CP-element group 282: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Update/ca
      -- CP-element group 282: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/Update/$exit
      -- 
    ca_3435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_986_inst_ack_1, ack => convolution3D_CP_1120_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	287 
    -- CP-element group 283:  members (5) 
      -- CP-element group 283: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_req
      -- CP-element group 283: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/$exit
      -- CP-element group 283: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/$exit
      -- CP-element group 283: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/$exit
      -- CP-element group 283: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_980/phi_stmt_980_sources/type_cast_986/SplitProtocol/$exit
      -- 
    phi_stmt_980_req_3436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_980_req_3436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(283), ack => phi_stmt_980_req_1); -- 
    convolution3D_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(281) & convolution3D_CP_1120_elements(282);
      gj_convolution3D_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	138 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Sample/ra
      -- CP-element group 284: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Sample/$exit
      -- 
    ra_3453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_993_inst_ack_0, ack => convolution3D_CP_1120_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	138 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Update/ca
      -- CP-element group 285: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/Update/$exit
      -- 
    ca_3458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_993_inst_ack_1, ack => convolution3D_CP_1120_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (5) 
      -- CP-element group 286: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/$exit
      -- CP-element group 286: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/$exit
      -- CP-element group 286: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_req
      -- CP-element group 286: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/SplitProtocol/$exit
      -- CP-element group 286: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_987/phi_stmt_987_sources/type_cast_993/$exit
      -- 
    phi_stmt_987_req_3459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_987_req_3459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(286), ack => phi_stmt_987_req_1); -- 
    convolution3D_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(284) & convolution3D_CP_1120_elements(285);
      gj_convolution3D_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	283 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (1) 
      -- CP-element group 287: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(283) & convolution3D_CP_1120_elements(286);
      gj_convolution3D_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  merge  fork  transition  place  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	280 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (2) 
      -- CP-element group 288: 	 branch_block_stmt_436/merge_stmt_979_PhiAck/$entry
      -- CP-element group 288: 	 branch_block_stmt_436/merge_stmt_979_PhiReqMerge
      -- 
    convolution3D_CP_1120_elements(288) <= OrReduce(convolution3D_CP_1120_elements(280) & convolution3D_CP_1120_elements(287));
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (1) 
      -- CP-element group 289: 	 branch_block_stmt_436/merge_stmt_979_PhiAck/phi_stmt_980_ack
      -- 
    phi_stmt_980_ack_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_980_ack_0, ack => convolution3D_CP_1120_elements(289)); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (1) 
      -- CP-element group 290: 	 branch_block_stmt_436/merge_stmt_979_PhiAck/phi_stmt_987_ack
      -- 
    phi_stmt_987_ack_3465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_987_ack_0, ack => convolution3D_CP_1120_elements(290)); -- 
    -- CP-element group 291:  join  fork  transition  place  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	131 
    -- CP-element group 291: 	134 
    -- CP-element group 291: 	135 
    -- CP-element group 291: 	136 
    -- CP-element group 291:  members (16) 
      -- CP-element group 291: 	 branch_block_stmt_436/merge_stmt_979__exit__
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033__entry__
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/$entry
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/RPIPE_maxpool_input_pipe_1008_Sample/rr
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_update_start_
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1012_Update/cr
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_update_start_
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Sample/rr
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1000_to_assign_stmt_1033/type_cast_1027_Update/cr
      -- CP-element group 291: 	 branch_block_stmt_436/merge_stmt_979_PhiAck/$exit
      -- 
    rr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(291), ack => RPIPE_maxpool_input_pipe_1008_inst_req_0); -- 
    cr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(291), ack => type_cast_1012_inst_req_1); -- 
    rr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(291), ack => type_cast_1027_inst_req_0); -- 
    cr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(291), ack => type_cast_1027_inst_req_1); -- 
    convolution3D_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(289) & convolution3D_CP_1120_elements(290);
      gj_convolution3D_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	139 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Sample/ra
      -- CP-element group 292: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Sample/$exit
      -- 
    ra_3489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1044_inst_ack_0, ack => convolution3D_CP_1120_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	139 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (2) 
      -- CP-element group 293: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/Update/ca
      -- 
    ca_3494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1044_inst_ack_1, ack => convolution3D_CP_1120_elements(293)); -- 
    -- CP-element group 294:  join  transition  place  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (8) 
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_req
      -- CP-element group 294: 	 branch_block_stmt_436/merge_stmt_1040_PhiAck/$entry
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/SplitProtocol/$exit
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1044/$exit
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/$exit
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1041/$exit
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 294: 	 branch_block_stmt_436/merge_stmt_1040_PhiReqMerge
      -- 
    phi_stmt_1041_req_3495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1041_req_3495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(294), ack => phi_stmt_1041_req_0); -- 
    convolution3D_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(292) & convolution3D_CP_1120_elements(293);
      gj_convolution3D_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	140 
    -- CP-element group 295: 	141 
    -- CP-element group 295: 	143 
    -- CP-element group 295: 	145 
    -- CP-element group 295:  members (29) 
      -- CP-element group 295: 	 branch_block_stmt_436/merge_stmt_1040__exit__
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079__entry__
      -- CP-element group 295: 	 branch_block_stmt_436/merge_stmt_1040_PhiAck/$exit
      -- CP-element group 295: 	 branch_block_stmt_436/merge_stmt_1040_PhiAck/phi_stmt_1041_ack
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_update_start_
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_resized_1
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_scaled_1
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_computed_1
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_resize_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_resize_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_resize_1/index_resize_req
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_resize_1/index_resize_ack
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_scale_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_scale_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_scale_1/scale_rename_req
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_index_scale_1/scale_rename_ack
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_update_start
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Sample/req
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/array_obj_ref_1073_final_index_sum_regn_Update/req
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/addr_of_1074_complete/req
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_update_start_
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/word_access_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/word_access_complete/word_0/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1079/ptr_deref_1077_Update/word_access_complete/word_0/cr
      -- 
    phi_stmt_1041_ack_3500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1041_ack_0, ack => convolution3D_CP_1120_elements(295)); -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(295), ack => array_obj_ref_1073_index_offset_req_0); -- 
    req_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(295), ack => array_obj_ref_1073_index_offset_req_1); -- 
    req_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(295), ack => addr_of_1074_final_reg_req_1); -- 
    cr_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(295), ack => ptr_deref_1077_store_0_req_1); -- 
    -- CP-element group 296:  merge  fork  transition  place  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	129 
    -- CP-element group 296: 	146 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	147 
    -- CP-element group 296: 	148 
    -- CP-element group 296: 	149 
    -- CP-element group 296: 	150 
    -- CP-element group 296: 	151 
    -- CP-element group 296: 	152 
    -- CP-element group 296: 	153 
    -- CP-element group 296: 	154 
    -- CP-element group 296:  members (31) 
      -- CP-element group 296: 	 branch_block_stmt_436/merge_stmt_1081__exit__
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133__entry__
      -- CP-element group 296: 	 branch_block_stmt_436/merge_stmt_1081_PhiAck/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/merge_stmt_1081_PhiAck/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/merge_stmt_1081_PhiAck/dummy
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_update_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Sample/rr
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Update/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1084_Update/cr
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_update_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Sample/rr
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Update/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1088_Update/cr
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_update_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Sample/rr
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Update/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1092_Update/cr
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_update_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Sample/rr
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Update/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1085_to_assign_stmt_1133/type_cast_1096_Update/cr
      -- CP-element group 296: 	 branch_block_stmt_436/merge_stmt_1081_PhiReqMerge
      -- 
    rr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1084_inst_req_0); -- 
    cr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1084_inst_req_1); -- 
    rr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1088_inst_req_0); -- 
    cr_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1088_inst_req_1); -- 
    rr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1092_inst_req_0); -- 
    cr_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1092_inst_req_1); -- 
    rr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1096_inst_req_0); -- 
    cr_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1096_inst_req_1); -- 
    convolution3D_CP_1120_elements(296) <= OrReduce(convolution3D_CP_1120_elements(129) & convolution3D_CP_1120_elements(146));
    -- CP-element group 297:  transition  output  delay-element  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	170 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	301 
    -- CP-element group 297:  members (5) 
      -- CP-element group 297: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- CP-element group 297: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1214/$exit
      -- CP-element group 297: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/$exit
      -- CP-element group 297: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1218_konst_delay_trans
      -- CP-element group 297: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_req
      -- 
    phi_stmt_1214_req_3534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1214_req_3534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(297), ack => phi_stmt_1214_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(297) is a control-delay.
    cp_element_297_delay: control_delay_element  generic map(name => " 297_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(170), ack => convolution3D_CP_1120_elements(297), clk => clk, reset =>reset);
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	212 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (2) 
      -- CP-element group 298: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Sample/$exit
      -- CP-element group 298: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Sample/ra
      -- 
    ra_3554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_0, ack => convolution3D_CP_1120_elements(298)); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	212 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (2) 
      -- CP-element group 299: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Update/$exit
      -- CP-element group 299: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/Update/ca
      -- 
    ca_3559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_1, ack => convolution3D_CP_1120_elements(299)); -- 
    -- CP-element group 300:  join  transition  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/SplitProtocol/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/type_cast_1220/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_sources/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1214/phi_stmt_1214_req
      -- 
    phi_stmt_1214_req_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1214_req_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(300), ack => phi_stmt_1214_req_1); -- 
    convolution3D_cp_element_group_300: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_300"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(298) & convolution3D_CP_1120_elements(299);
      gj_convolution3D_cp_element_group_300 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(300), clk => clk, reset => reset); --
    end block;
    -- CP-element group 301:  merge  transition  place  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	297 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (2) 
      -- CP-element group 301: 	 branch_block_stmt_436/merge_stmt_1213_PhiReqMerge
      -- CP-element group 301: 	 branch_block_stmt_436/merge_stmt_1213_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(301) <= OrReduce(convolution3D_CP_1120_elements(297) & convolution3D_CP_1120_elements(300));
    -- CP-element group 302:  fork  transition  place  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	171 
    -- CP-element group 302: 	172 
    -- CP-element group 302: 	174 
    -- CP-element group 302: 	175 
    -- CP-element group 302: 	178 
    -- CP-element group 302: 	182 
    -- CP-element group 302: 	186 
    -- CP-element group 302: 	190 
    -- CP-element group 302: 	194 
    -- CP-element group 302: 	198 
    -- CP-element group 302: 	202 
    -- CP-element group 302: 	206 
    -- CP-element group 302: 	209 
    -- CP-element group 302:  members (56) 
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_scale_1/scale_rename_ack
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_scale_1/$exit
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_resize_1/index_resize_ack
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_scale_1/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_scale_1/scale_rename_req
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1265_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1234_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_update_start
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Update/req
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/merge_stmt_1213__exit__
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376__entry__
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_resize_1/index_resize_req
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_resize_1/$exit
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_resize_1/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1283_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1319_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/RPIPE_maxpool_input_pipe_1230_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1247_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_final_index_sum_regn_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_complete/req
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1301_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/addr_of_1227_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_resized_1
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_scaled_1
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/array_obj_ref_1226_index_computed_1
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1337_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/type_cast_1355_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_update_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/word_access_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/word_access_complete/word_0/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1228_to_assign_stmt_1376/ptr_deref_1363_Update/word_access_complete/word_0/cr
      -- CP-element group 302: 	 branch_block_stmt_436/merge_stmt_1213_PhiAck/phi_stmt_1214_ack
      -- CP-element group 302: 	 branch_block_stmt_436/merge_stmt_1213_PhiAck/$exit
      -- 
    phi_stmt_1214_ack_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1214_ack_0, ack => convolution3D_CP_1120_elements(302)); -- 
    cr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1265_inst_req_1); -- 
    cr_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1234_inst_req_1); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => array_obj_ref_1226_index_offset_req_1); -- 
    cr_2654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1283_inst_req_1); -- 
    rr_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => RPIPE_maxpool_input_pipe_1230_inst_req_0); -- 
    cr_2598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1247_inst_req_1); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1319_inst_req_1); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => array_obj_ref_1226_index_offset_req_0); -- 
    req_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => addr_of_1227_final_reg_req_1); -- 
    cr_2682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1301_inst_req_1); -- 
    cr_2738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1337_inst_req_1); -- 
    cr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => type_cast_1355_inst_req_1); -- 
    cr_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => ptr_deref_1363_store_0_req_1); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	211 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	305 
    -- CP-element group 303:  members (2) 
      -- CP-element group 303: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Sample/ra
      -- CP-element group 303: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Sample/$exit
      -- 
    ra_3597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_0, ack => convolution3D_CP_1120_elements(303)); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	211 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (2) 
      -- CP-element group 304: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Update/ca
      -- CP-element group 304: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/Update/$exit
      -- 
    ca_3602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_1, ack => convolution3D_CP_1120_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	303 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_req
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/SplitProtocol/$exit
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1411/$exit
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$exit
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1408/$exit
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- 
    phi_stmt_1408_req_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1408_req_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(305), ack => phi_stmt_1408_req_0); -- 
    convolution3D_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(303) & convolution3D_CP_1120_elements(304);
      gj_convolution3D_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  transition  output  delay-element  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	157 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (5) 
      -- CP-element group 306: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414_konst_delay_trans
      -- CP-element group 306: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_req
      -- CP-element group 306: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$exit
      -- CP-element group 306: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1408/$exit
      -- CP-element group 306: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/$exit
      -- 
    phi_stmt_1408_req_3614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1408_req_3614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(306), ack => phi_stmt_1408_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(306) is a control-delay.
    cp_element_306_delay: control_delay_element  generic map(name => " 306_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(157), ack => convolution3D_CP_1120_elements(306), clk => clk, reset =>reset);
    -- CP-element group 307:  merge  transition  place  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (2) 
      -- CP-element group 307: 	 branch_block_stmt_436/merge_stmt_1407_PhiReqMerge
      -- CP-element group 307: 	 branch_block_stmt_436/merge_stmt_1407_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(307) <= OrReduce(convolution3D_CP_1120_elements(305) & convolution3D_CP_1120_elements(306));
    -- CP-element group 308:  branch  transition  place  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	213 
    -- CP-element group 308: 	214 
    -- CP-element group 308:  members (15) 
      -- CP-element group 308: 	 branch_block_stmt_436/R_tobool218_1429_place
      -- CP-element group 308: 	 branch_block_stmt_436/merge_stmt_1407__exit__
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1421_to_assign_stmt_1427__entry__
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1421_to_assign_stmt_1427__exit__
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1428__entry__
      -- CP-element group 308: 	 branch_block_stmt_436/merge_stmt_1407_PhiAck/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/merge_stmt_1407_PhiAck/phi_stmt_1408_ack
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1421_to_assign_stmt_1427/$entry
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1421_to_assign_stmt_1427/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1428_dead_link/$entry
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1428_eval_test/$entry
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1428_eval_test/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1428_eval_test/branch_req
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1428_if_link/$entry
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1428_else_link/$entry
      -- 
    phi_stmt_1408_ack_3619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1408_ack_0, ack => convolution3D_CP_1120_elements(308)); -- 
    branch_req_2850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(308), ack => if_stmt_1428_branch_req_0); -- 
    -- CP-element group 309:  transition  output  delay-element  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	216 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (4) 
      -- CP-element group 309: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_req
      -- CP-element group 309: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1457_konst_delay_trans
      -- CP-element group 309: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/$exit
      -- CP-element group 309: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/$exit
      -- 
    phi_stmt_1453_req_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1453_req_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(309), ack => phi_stmt_1453_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(309) is a control-delay.
    cp_element_309_delay: control_delay_element  generic map(name => " 309_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(216), ack => convolution3D_CP_1120_elements(309), clk => clk, reset =>reset);
    -- CP-element group 310:  transition  output  delay-element  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	216 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (4) 
      -- CP-element group 310: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_req
      -- CP-element group 310: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1464_konst_delay_trans
      -- CP-element group 310: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/$exit
      -- CP-element group 310: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/$exit
      -- 
    phi_stmt_1460_req_3650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1460_req_3650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(310), ack => phi_stmt_1460_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(310) is a control-delay.
    cp_element_310_delay: control_delay_element  generic map(name => " 310_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(216), ack => convolution3D_CP_1120_elements(310), clk => clk, reset =>reset);
    -- CP-element group 311:  join  transition  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	319 
    -- CP-element group 311:  members (1) 
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(309) & convolution3D_CP_1120_elements(310);
      gj_convolution3D_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	224 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (2) 
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Sample/ra
      -- 
    ra_3670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1459_inst_ack_0, ack => convolution3D_CP_1120_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	224 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (2) 
      -- CP-element group 313: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/Update/ca
      -- 
    ca_3675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1459_inst_ack_1, ack => convolution3D_CP_1120_elements(313)); -- 
    -- CP-element group 314:  join  transition  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	318 
    -- CP-element group 314:  members (5) 
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/SplitProtocol/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/type_cast_1459/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_sources/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1453/phi_stmt_1453_req
      -- 
    phi_stmt_1453_req_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1453_req_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(314), ack => phi_stmt_1453_req_1); -- 
    convolution3D_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(312) & convolution3D_CP_1120_elements(313);
      gj_convolution3D_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	224 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Sample/ra
      -- CP-element group 315: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Sample/$exit
      -- 
    ra_3693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_0, ack => convolution3D_CP_1120_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	224 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/Update/ca
      -- 
    ca_3698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_1, ack => convolution3D_CP_1120_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (5) 
      -- CP-element group 317: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/$exit
      -- CP-element group 317: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/$exit
      -- CP-element group 317: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/$exit
      -- CP-element group 317: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_sources/type_cast_1466/SplitProtocol/$exit
      -- CP-element group 317: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1460/phi_stmt_1460_req
      -- 
    phi_stmt_1460_req_3699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1460_req_3699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(317), ack => phi_stmt_1460_req_1); -- 
    convolution3D_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(315) & convolution3D_CP_1120_elements(316);
      gj_convolution3D_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  transition  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	314 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (1) 
      -- CP-element group 318: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(314) & convolution3D_CP_1120_elements(317);
      gj_convolution3D_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  merge  fork  transition  place  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	311 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_436/merge_stmt_1452_PhiReqMerge
      -- CP-element group 319: 	 branch_block_stmt_436/merge_stmt_1452_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(319) <= OrReduce(convolution3D_CP_1120_elements(311) & convolution3D_CP_1120_elements(318));
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	322 
    -- CP-element group 320:  members (1) 
      -- CP-element group 320: 	 branch_block_stmt_436/merge_stmt_1452_PhiAck/phi_stmt_1453_ack
      -- 
    phi_stmt_1453_ack_3704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1453_ack_0, ack => convolution3D_CP_1120_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (1) 
      -- CP-element group 321: 	 branch_block_stmt_436/merge_stmt_1452_PhiAck/phi_stmt_1460_ack
      -- 
    phi_stmt_1460_ack_3705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1460_ack_0, ack => convolution3D_CP_1120_elements(321)); -- 
    -- CP-element group 322:  join  fork  transition  place  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	320 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	217 
    -- CP-element group 322: 	220 
    -- CP-element group 322: 	221 
    -- CP-element group 322: 	222 
    -- CP-element group 322:  members (16) 
      -- CP-element group 322: 	 branch_block_stmt_436/merge_stmt_1452__exit__
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506__entry__
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/RPIPE_maxpool_input_pipe_1481_Sample/rr
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_update_start_
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1485_Update/cr
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_update_start_
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Sample/rr
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1473_to_assign_stmt_1506/type_cast_1500_Update/cr
      -- CP-element group 322: 	 branch_block_stmt_436/merge_stmt_1452_PhiAck/$exit
      -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(322), ack => RPIPE_maxpool_input_pipe_1481_inst_req_0); -- 
    cr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(322), ack => type_cast_1485_inst_req_1); -- 
    rr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(322), ack => type_cast_1500_inst_req_0); -- 
    cr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(322), ack => type_cast_1500_inst_req_1); -- 
    convolution3D_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(320) & convolution3D_CP_1120_elements(321);
      gj_convolution3D_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	225 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (2) 
      -- CP-element group 323: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Sample/ra
      -- 
    ra_3729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1517_inst_ack_0, ack => convolution3D_CP_1120_elements(323)); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	225 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (2) 
      -- CP-element group 324: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Update/ca
      -- CP-element group 324: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/Update/$exit
      -- 
    ca_3734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1517_inst_ack_1, ack => convolution3D_CP_1120_elements(324)); -- 
    -- CP-element group 325:  join  transition  place  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (8) 
      -- CP-element group 325: 	 branch_block_stmt_436/merge_stmt_1513_PhiReqMerge
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/SplitProtocol/$exit
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/type_cast_1517/$exit
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_sources/$exit
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/$exit
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/$exit
      -- CP-element group 325: 	 branch_block_stmt_436/merge_stmt_1513_PhiAck/$entry
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1514/phi_stmt_1514_req
      -- 
    phi_stmt_1514_req_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1514_req_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(325), ack => phi_stmt_1514_req_0); -- 
    convolution3D_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(323) & convolution3D_CP_1120_elements(324);
      gj_convolution3D_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	226 
    -- CP-element group 326: 	227 
    -- CP-element group 326: 	229 
    -- CP-element group 326: 	231 
    -- CP-element group 326:  members (29) 
      -- CP-element group 326: 	 branch_block_stmt_436/merge_stmt_1513__exit__
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552__entry__
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_update_start_
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_resized_1
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_scaled_1
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_computed_1
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_resize_1/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_resize_1/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_resize_1/index_resize_req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_resize_1/index_resize_ack
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_scale_1/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_scale_1/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_scale_1/scale_rename_req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_index_scale_1/scale_rename_ack
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_update_start
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Sample/req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/array_obj_ref_1546_final_index_sum_regn_Update/req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_complete/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/addr_of_1547_complete/req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_update_start_
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/word_access_complete/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/word_access_complete/word_0/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1524_to_assign_stmt_1552/ptr_deref_1550_Update/word_access_complete/word_0/cr
      -- CP-element group 326: 	 branch_block_stmt_436/merge_stmt_1513_PhiAck/phi_stmt_1514_ack
      -- CP-element group 326: 	 branch_block_stmt_436/merge_stmt_1513_PhiAck/$exit
      -- 
    phi_stmt_1514_ack_3740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1514_ack_0, ack => convolution3D_CP_1120_elements(326)); -- 
    req_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => array_obj_ref_1546_index_offset_req_0); -- 
    req_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => array_obj_ref_1546_index_offset_req_1); -- 
    req_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => addr_of_1547_final_reg_req_1); -- 
    cr_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => ptr_deref_1550_store_0_req_1); -- 
    -- CP-element group 327:  merge  fork  transition  place  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	213 
    -- CP-element group 327: 	232 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	233 
    -- CP-element group 327: 	234 
    -- CP-element group 327:  members (13) 
      -- CP-element group 327: 	 branch_block_stmt_436/merge_stmt_1554__exit__
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557__entry__
      -- CP-element group 327: 	 branch_block_stmt_436/merge_stmt_1554_PhiReqMerge
      -- CP-element group 327: 	 branch_block_stmt_436/merge_stmt_1554_PhiAck/dummy
      -- CP-element group 327: 	 branch_block_stmt_436/merge_stmt_1554_PhiAck/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/merge_stmt_1554_PhiAck/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_sample_start_
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_update_start_
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Sample/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Sample/crr
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/call_stmt_1557/call_stmt_1557_Update/ccr
      -- 
    crr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(327), ack => call_stmt_1557_call_req_0); -- 
    ccr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(327), ack => call_stmt_1557_call_req_1); -- 
    convolution3D_CP_1120_elements(327) <= OrReduce(convolution3D_CP_1120_elements(213) & convolution3D_CP_1120_elements(232));
    -- CP-element group 328:  transition  output  delay-element  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	245 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	332 
    -- CP-element group 328:  members (5) 
      -- CP-element group 328: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$exit
      -- CP-element group 328: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1630_konst_delay_trans
      -- CP-element group 328: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_req
      -- CP-element group 328: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1624/$exit
      -- CP-element group 328: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1624_req_3762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1624_req_3762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(328), ack => phi_stmt_1624_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(328) is a control-delay.
    cp_element_328_delay: control_delay_element  generic map(name => " 328_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(245), ack => convolution3D_CP_1120_elements(328), clk => clk, reset =>reset);
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	257 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (2) 
      -- CP-element group 329: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/ra
      -- CP-element group 329: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/$exit
      -- 
    ra_3782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_0, ack => convolution3D_CP_1120_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	257 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (2) 
      -- CP-element group 330: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/ca
      -- CP-element group 330: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/$exit
      -- 
    ca_3787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_1, ack => convolution3D_CP_1120_elements(330)); -- 
    -- CP-element group 331:  join  transition  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_req
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$exit
      -- 
    phi_stmt_1624_req_3788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1624_req_3788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => phi_stmt_1624_req_0); -- 
    convolution3D_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(329) & convolution3D_CP_1120_elements(330);
      gj_convolution3D_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  merge  transition  place  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	328 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_436/merge_stmt_1623_PhiReqMerge
      -- CP-element group 332: 	 branch_block_stmt_436/merge_stmt_1623_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(332) <= OrReduce(convolution3D_CP_1120_elements(328) & convolution3D_CP_1120_elements(331));
    -- CP-element group 333:  fork  transition  place  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	246 
    -- CP-element group 333: 	247 
    -- CP-element group 333: 	248 
    -- CP-element group 333: 	249 
    -- CP-element group 333: 	252 
    -- CP-element group 333: 	253 
    -- CP-element group 333: 	254 
    -- CP-element group 333:  members (26) 
      -- CP-element group 333: 	 branch_block_stmt_436/merge_stmt_1623_PhiAck/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/merge_stmt_1623__exit__
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670__entry__
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_update_start_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Sample/rr
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1644_Update/cr
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_update_start_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Sample/rr
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/type_cast_1648_Update/cr
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_update_start_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1652_Update/ccr
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_update_start_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Sample/crr
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1636_to_assign_stmt_1670/call_stmt_1659_Update/ccr
      -- CP-element group 333: 	 branch_block_stmt_436/merge_stmt_1623_PhiAck/phi_stmt_1624_ack
      -- 
    phi_stmt_1624_ack_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1624_ack_0, ack => convolution3D_CP_1120_elements(333)); -- 
    rr_3142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => type_cast_1644_inst_req_0); -- 
    cr_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => type_cast_1644_inst_req_1); -- 
    rr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => type_cast_1648_inst_req_0); -- 
    cr_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => type_cast_1648_inst_req_1); -- 
    ccr_3175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => call_stmt_1652_call_req_1); -- 
    crr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => call_stmt_1659_call_req_0); -- 
    ccr_3189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => call_stmt_1659_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1125_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1403_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_934_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1051 : std_logic_vector(63 downto 0);
    signal R_indvar350_1225_resized : std_logic_vector(13 downto 0);
    signal R_indvar350_1225_scaled : std_logic_vector(13 downto 0);
    signal R_indvar364_756_resized : std_logic_vector(13 downto 0);
    signal R_indvar364_756_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1072_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1072_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1545_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1545_scaled : std_logic_vector(13 downto 0);
    signal add102_802 : std_logic_vector(63 downto 0);
    signal add108_820 : std_logic_vector(63 downto 0);
    signal add114_838 : std_logic_vector(63 downto 0);
    signal add120_856 : std_logic_vector(63 downto 0);
    signal add1216x_xi308_1530 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1057 : std_logic_vector(63 downto 0);
    signal add126_874 : std_logic_vector(63 downto 0);
    signal add132_892 : std_logic_vector(63 downto 0);
    signal add13_486 : std_logic_vector(15 downto 0);
    signal add171_1253 : std_logic_vector(63 downto 0);
    signal add177_1271 : std_logic_vector(63 downto 0);
    signal add183_1289 : std_logic_vector(63 downto 0);
    signal add189_1307 : std_logic_vector(63 downto 0);
    signal add195_1325 : std_logic_vector(63 downto 0);
    signal add201_1343 : std_logic_vector(63 downto 0);
    signal add207_1361 : std_logic_vector(63 downto 0);
    signal add23_511 : std_logic_vector(15 downto 0);
    signal add33_536 : std_logic_vector(15 downto 0);
    signal add43_561 : std_logic_vector(15 downto 0);
    signal add53_586 : std_logic_vector(15 downto 0);
    signal add63_611 : std_logic_vector(15 downto 0);
    signal add73_636 : std_logic_vector(15 downto 0);
    signal add96_784 : std_logic_vector(63 downto 0);
    signal add_461 : std_logic_vector(31 downto 0);
    signal addx_xi299_1491 : std_logic_vector(63 downto 0);
    signal addx_xi_1018 : std_logic_vector(63 downto 0);
    signal and217_1421 : std_logic_vector(63 downto 0);
    signal and_952 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1073_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1073_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1073_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1073_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1073_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1073_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1226_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1226_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1226_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1226_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1226_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1226_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1546_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1546_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1546_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1546_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1546_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1546_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_757_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_757_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_757_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_757_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_757_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_757_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1075 : std_logic_vector(31 downto 0);
    signal arrayidx211_1228 : std_logic_vector(31 downto 0);
    signal arrayidx226_1548 : std_logic_vector(31 downto 0);
    signal arrayidx_759 : std_logic_vector(31 downto 0);
    signal call105_811 : std_logic_vector(7 downto 0);
    signal call111_829 : std_logic_vector(7 downto 0);
    signal call117_847 : std_logic_vector(7 downto 0);
    signal call11_477 : std_logic_vector(7 downto 0);
    signal call123_865 : std_logic_vector(7 downto 0);
    signal call129_883 : std_logic_vector(7 downto 0);
    signal call164_1231 : std_logic_vector(7 downto 0);
    signal call168_1244 : std_logic_vector(7 downto 0);
    signal call16_489 : std_logic_vector(7 downto 0);
    signal call174_1262 : std_logic_vector(7 downto 0);
    signal call180_1280 : std_logic_vector(7 downto 0);
    signal call186_1298 : std_logic_vector(7 downto 0);
    signal call192_1316 : std_logic_vector(7 downto 0);
    signal call198_1334 : std_logic_vector(7 downto 0);
    signal call204_1352 : std_logic_vector(7 downto 0);
    signal call21_502 : std_logic_vector(7 downto 0);
    signal call229_1557 : std_logic_vector(63 downto 0);
    signal call26_514 : std_logic_vector(7 downto 0);
    signal call284_1685 : std_logic_vector(63 downto 0);
    signal call2_452 : std_logic_vector(7 downto 0);
    signal call31_527 : std_logic_vector(7 downto 0);
    signal call36_539 : std_logic_vector(7 downto 0);
    signal call41_552 : std_logic_vector(7 downto 0);
    signal call46_564 : std_logic_vector(7 downto 0);
    signal call51_577 : std_logic_vector(7 downto 0);
    signal call56_589 : std_logic_vector(7 downto 0);
    signal call61_602 : std_logic_vector(7 downto 0);
    signal call66_614 : std_logic_vector(7 downto 0);
    signal call6_464 : std_logic_vector(7 downto 0);
    signal call71_627 : std_logic_vector(7 downto 0);
    signal call89_762 : std_logic_vector(7 downto 0);
    signal call93_775 : std_logic_vector(7 downto 0);
    signal call99_793 : std_logic_vector(7 downto 0);
    signal call_439 : std_logic_vector(7 downto 0);
    signal callx_xi297_1482 : std_logic_vector(7 downto 0);
    signal callx_xi_1009 : std_logic_vector(7 downto 0);
    signal cmp161317_1133 : std_logic_vector(0 downto 0);
    signal cmp321_666 : std_logic_vector(0 downto 0);
    signal cmpx_xi302_1506 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1033 : std_logic_vector(0 downto 0);
    signal conv101_797 : std_logic_vector(63 downto 0);
    signal conv107_815 : std_logic_vector(63 downto 0);
    signal conv113_833 : std_logic_vector(63 downto 0);
    signal conv119_851 : std_logic_vector(63 downto 0);
    signal conv125_869 : std_logic_vector(63 downto 0);
    signal conv12_481 : std_logic_vector(15 downto 0);
    signal conv131_887 : std_logic_vector(63 downto 0);
    signal conv145_1085 : std_logic_vector(63 downto 0);
    signal conv147_1089 : std_logic_vector(63 downto 0);
    signal conv150_1093 : std_logic_vector(63 downto 0);
    signal conv153_1097 : std_logic_vector(63 downto 0);
    signal conv155_1127 : std_logic_vector(63 downto 0);
    signal conv165_1235 : std_logic_vector(63 downto 0);
    signal conv170_1248 : std_logic_vector(63 downto 0);
    signal conv176_1266 : std_logic_vector(63 downto 0);
    signal conv182_1284 : std_logic_vector(63 downto 0);
    signal conv188_1302 : std_logic_vector(63 downto 0);
    signal conv194_1320 : std_logic_vector(63 downto 0);
    signal conv19_493 : std_logic_vector(15 downto 0);
    signal conv1_443 : std_logic_vector(31 downto 0);
    signal conv200_1338 : std_logic_vector(63 downto 0);
    signal conv206_1356 : std_logic_vector(63 downto 0);
    signal conv22_506 : std_logic_vector(15 downto 0);
    signal conv230_1682 : std_logic_vector(63 downto 0);
    signal conv255_1645 : std_logic_vector(63 downto 0);
    signal conv261_1649 : std_logic_vector(63 downto 0);
    signal conv285_1690 : std_logic_vector(63 downto 0);
    signal conv29_518 : std_logic_vector(15 downto 0);
    signal conv2x_xi292_1444 : std_logic_vector(31 downto 0);
    signal conv2x_xi_971 : std_logic_vector(31 downto 0);
    signal conv32_531 : std_logic_vector(15 downto 0);
    signal conv39_543 : std_logic_vector(15 downto 0);
    signal conv3_456 : std_logic_vector(31 downto 0);
    signal conv42_556 : std_logic_vector(15 downto 0);
    signal conv49_568 : std_logic_vector(15 downto 0);
    signal conv52_581 : std_logic_vector(15 downto 0);
    signal conv59_593 : std_logic_vector(15 downto 0);
    signal conv5x_xi298_1486 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1013 : std_logic_vector(63 downto 0);
    signal conv62_606 : std_logic_vector(15 downto 0);
    signal conv69_618 : std_logic_vector(15 downto 0);
    signal conv72_631 : std_logic_vector(15 downto 0);
    signal conv79_640 : std_logic_vector(31 downto 0);
    signal conv81_644 : std_logic_vector(31 downto 0);
    signal conv83_660 : std_logic_vector(63 downto 0);
    signal conv90_766 : std_logic_vector(63 downto 0);
    signal conv95_779 : std_logic_vector(63 downto 0);
    signal conv9_468 : std_logic_vector(15 downto 0);
    signal convx_xi301_1501 : std_logic_vector(31 downto 0);
    signal convx_xi_1028 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi296_1460 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_987 : std_logic_vector(63 downto 0);
    signal exitcond32_907 : std_logic_vector(0 downto 0);
    signal exitcond5_1670 : std_logic_vector(0 downto 0);
    signal exitcond_1376 : std_logic_vector(0 downto 0);
    signal iNsTr_34_1006 : std_logic_vector(15 downto 0);
    signal iNsTr_54_1440 : std_logic_vector(63 downto 0);
    signal iNsTr_62_1479 : std_logic_vector(15 downto 0);
    signal iNsTr_70_1524 : std_logic_vector(63 downto 0);
    signal indvar350_1214 : std_logic_vector(63 downto 0);
    signal indvar364_745 : std_logic_vector(63 downto 0);
    signal indvar_1624 : std_logic_vector(31 downto 0);
    signal indvarx_xnext351_1371 : std_logic_vector(63 downto 0);
    signal indvarx_xnext365_902 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1665 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_939 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1408 : std_logic_vector(63 downto 0);
    signal mul148_1102 : std_logic_vector(63 downto 0);
    signal mul151_1107 : std_logic_vector(63 downto 0);
    signal mul154_1112 : std_logic_vector(63 downto 0);
    signal mul236_1563 : std_logic_vector(15 downto 0);
    signal mul249_1568 : std_logic_vector(15 downto 0);
    signal mul254_1636 : std_logic_vector(31 downto 0);
    signal mul260_1641 : std_logic_vector(31 downto 0);
    signal mul82_654 : std_logic_vector(31 downto 0);
    signal mul_649 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi295_1453 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_980 : std_logic_vector(15 downto 0);
    signal phitmp325_1405 : std_logic_vector(63 downto 0);
    signal phitmp_936 : std_logic_vector(63 downto 0);
    signal ptr_deref_1077_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1077_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1077_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1077_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1077_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1077_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1363_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1363_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1363_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1363_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1363_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1363_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1550_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1550_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1550_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1550_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1550_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1550_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_894_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_894_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_894_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_894_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_894_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_894_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1118 : std_logic_vector(63 downto 0);
    signal sh_promx_xi309_1536 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1063 : std_logic_vector(63 downto 0);
    signal shl104_808 : std_logic_vector(63 downto 0);
    signal shl10_474 : std_logic_vector(15 downto 0);
    signal shl110_826 : std_logic_vector(63 downto 0);
    signal shl116_844 : std_logic_vector(63 downto 0);
    signal shl122_862 : std_logic_vector(63 downto 0);
    signal shl128_880 : std_logic_vector(63 downto 0);
    signal shl14x_xi310_1541 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1068 : std_logic_vector(63 downto 0);
    signal shl167_1241 : std_logic_vector(63 downto 0);
    signal shl173_1259 : std_logic_vector(63 downto 0);
    signal shl179_1277 : std_logic_vector(63 downto 0);
    signal shl185_1295 : std_logic_vector(63 downto 0);
    signal shl191_1313 : std_logic_vector(63 downto 0);
    signal shl197_1331 : std_logic_vector(63 downto 0);
    signal shl203_1349 : std_logic_vector(63 downto 0);
    signal shl20_499 : std_logic_vector(15 downto 0);
    signal shl30_524 : std_logic_vector(15 downto 0);
    signal shl40_549 : std_logic_vector(15 downto 0);
    signal shl50_574 : std_logic_vector(15 downto 0);
    signal shl60_599 : std_logic_vector(15 downto 0);
    signal shl70_624 : std_logic_vector(15 downto 0);
    signal shl8x_xi300_1497 : std_logic_vector(63 downto 0);
    signal shl8x_xi300x_xlcssa_1514 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1024 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1041 : std_logic_vector(63 downto 0);
    signal shl92_772 : std_logic_vector(63 downto 0);
    signal shl98_790 : std_logic_vector(63 downto 0);
    signal shl_449 : std_logic_vector(31 downto 0);
    signal shlx_xi293_1450 : std_logic_vector(31 downto 0);
    signal shlx_xi_977 : std_logic_vector(31 downto 0);
    signal sub269_1587 : std_logic_vector(15 downto 0);
    signal sub289_1695 : std_logic_vector(63 downto 0);
    signal sub_1581 : std_logic_vector(15 downto 0);
    signal tmp12_1156 : std_logic_vector(63 downto 0);
    signal tmp13_1160 : std_logic_vector(63 downto 0);
    signal tmp14_1165 : std_logic_vector(63 downto 0);
    signal tmp15_1169 : std_logic_vector(63 downto 0);
    signal tmp16_1174 : std_logic_vector(63 downto 0);
    signal tmp17_1178 : std_logic_vector(63 downto 0);
    signal tmp18_1183 : std_logic_vector(63 downto 0);
    signal tmp19_1187 : std_logic_vector(31 downto 0);
    signal tmp20_1192 : std_logic_vector(63 downto 0);
    signal tmp21_1198 : std_logic_vector(63 downto 0);
    signal tmp22_1204 : std_logic_vector(0 downto 0);
    signal tmp24_704 : std_logic_vector(31 downto 0);
    signal tmp25_709 : std_logic_vector(31 downto 0);
    signal tmp26_713 : std_logic_vector(31 downto 0);
    signal tmp27_718 : std_logic_vector(31 downto 0);
    signal tmp28_723 : std_logic_vector(63 downto 0);
    signal tmp29_729 : std_logic_vector(63 downto 0);
    signal tmp30_735 : std_logic_vector(0 downto 0);
    signal tmp326_1473 : std_logic_vector(15 downto 0);
    signal tmp327_1593 : std_logic_vector(15 downto 0);
    signal tmp345_1146 : std_logic_vector(63 downto 0);
    signal tmp346_1152 : std_logic_vector(0 downto 0);
    signal tmp347_1396 : std_logic_vector(63 downto 0);
    signal tmp354_678 : std_logic_vector(31 downto 0);
    signal tmp356_683 : std_logic_vector(31 downto 0);
    signal tmp357_688 : std_logic_vector(63 downto 0);
    signal tmp358_694 : std_logic_vector(63 downto 0);
    signal tmp359_700 : std_logic_vector(0 downto 0);
    signal tmp361_927 : std_logic_vector(63 downto 0);
    signal tmp3_1597 : std_logic_vector(31 downto 0);
    signal tmp4_1603 : std_logic_vector(31 downto 0);
    signal tmp6_1607 : std_logic_vector(31 downto 0);
    signal tmp7_1612 : std_logic_vector(15 downto 0);
    signal tmp8_1616 : std_logic_vector(31 downto 0);
    signal tmp9_1621 : std_logic_vector(31 downto 0);
    signal tmp_1000 : std_logic_vector(15 downto 0);
    signal tobool218_1427 : std_logic_vector(0 downto 0);
    signal tobool_958 : std_logic_vector(0 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1022_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1044_wire : std_logic_vector(63 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1055_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1061_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1121_wire : std_logic_vector(63 downto 0);
    signal type_cast_1124_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1131_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1150_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1190_wire : std_logic_vector(63 downto 0);
    signal type_cast_1196_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1202_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1209_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1218_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1220_wire : std_logic_vector(63 downto 0);
    signal type_cast_1239_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1257_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1275_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1293_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1311_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1329_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1347_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1369_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1388_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1394_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1399_wire : std_logic_vector(63 downto 0);
    signal type_cast_1402_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1411_wire : std_logic_vector(63 downto 0);
    signal type_cast_1414_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1419_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1425_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1448_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1457_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1459_wire : std_logic_vector(15 downto 0);
    signal type_cast_1464_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1466_wire : std_logic_vector(63 downto 0);
    signal type_cast_1471_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1477_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1495_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1517_wire : std_logic_vector(63 downto 0);
    signal type_cast_1522_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1528_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1534_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1574_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1579_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1585_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1591_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1601_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1627_wire : std_logic_vector(31 downto 0);
    signal type_cast_1630_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1663_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1680_wire : std_logic_vector(63 downto 0);
    signal type_cast_1688_wire : std_logic_vector(63 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_472_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_497_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_522_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_547_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_572_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_597_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_622_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_658_wire : std_logic_vector(63 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_686_wire : std_logic_vector(63 downto 0);
    signal type_cast_692_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_721_wire : std_logic_vector(63 downto 0);
    signal type_cast_727_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_733_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_740_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_749_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_751_wire : std_logic_vector(63 downto 0);
    signal type_cast_770_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_806_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_842_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_860_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_900_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_919_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_925_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_930_wire : std_logic_vector(63 downto 0);
    signal type_cast_933_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_942_wire : std_logic_vector(63 downto 0);
    signal type_cast_945_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_950_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_956_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_969_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_975_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_984_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_986_wire : std_logic_vector(15 downto 0);
    signal type_cast_991_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_993_wire : std_logic_vector(63 downto 0);
    signal type_cast_998_wire_constant : std_logic_vector(15 downto 0);
    signal umax23_1211 : std_logic_vector(63 downto 0);
    signal umax31_742 : std_logic_vector(63 downto 0);
    signal umax360_921 : std_logic_vector(63 downto 0);
    signal umax_1390 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1073_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1073_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1073_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1073_resized_base_address <= "00000000000000";
    array_obj_ref_1226_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1226_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1226_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1226_resized_base_address <= "00000000000000";
    array_obj_ref_1546_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1546_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1546_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1546_resized_base_address <= "00000000000000";
    array_obj_ref_757_constant_part_of_offset <= "00000000000000";
    array_obj_ref_757_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_757_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_757_resized_base_address <= "00000000000000";
    ptr_deref_1077_word_offset_0 <= "00000000000000";
    ptr_deref_1363_word_offset_0 <= "00000000000000";
    ptr_deref_1550_word_offset_0 <= "00000000000000";
    ptr_deref_894_word_offset_0 <= "00000000000000";
    type_cast_1004_wire_constant <= "0000000000000001";
    type_cast_1022_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1049_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1055_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1061_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1116_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1124_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1131_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1144_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1150_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1196_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1202_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1209_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1218_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1239_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1257_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1275_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1293_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1311_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1329_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1347_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1369_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1388_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1394_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1402_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1414_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1419_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1425_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1448_wire_constant <= "00000000000000000000000000000110";
    type_cast_1457_wire_constant <= "0000000000000000";
    type_cast_1464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1471_wire_constant <= "0000000000000001";
    type_cast_1477_wire_constant <= "0000000000000001";
    type_cast_1495_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1522_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1528_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1534_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1574_wire_constant <= "00101100";
    type_cast_1579_wire_constant <= "1111111111111111";
    type_cast_1585_wire_constant <= "1111111111111111";
    type_cast_1591_wire_constant <= "1111111111111111";
    type_cast_1601_wire_constant <= "00000000000000000000000000000001";
    type_cast_1630_wire_constant <= "00000000000000000000000000000000";
    type_cast_1663_wire_constant <= "00000000000000000000000000000001";
    type_cast_447_wire_constant <= "00000000000000000000000000001000";
    type_cast_472_wire_constant <= "0000000000001000";
    type_cast_497_wire_constant <= "0000000000001000";
    type_cast_522_wire_constant <= "0000000000001000";
    type_cast_547_wire_constant <= "0000000000001000";
    type_cast_572_wire_constant <= "0000000000001000";
    type_cast_597_wire_constant <= "0000000000001000";
    type_cast_622_wire_constant <= "0000000000001000";
    type_cast_664_wire_constant <= "00000000000000000000000000000011";
    type_cast_692_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_698_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_727_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_733_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_740_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_749_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_770_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_788_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_806_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_824_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_842_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_860_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_878_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_900_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_919_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_925_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_933_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_945_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_950_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_956_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_969_wire_constant <= "00000000000000000000000000000001";
    type_cast_975_wire_constant <= "00000000000000000000000000000110";
    type_cast_984_wire_constant <= "0000000000000000";
    type_cast_991_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_998_wire_constant <= "0000000000000001";
    phi_stmt_1041: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1044_wire;
      req(0) <= phi_stmt_1041_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1041",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1041_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1041,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1041
    phi_stmt_1214: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1218_wire_constant & type_cast_1220_wire;
      req <= phi_stmt_1214_req_0 & phi_stmt_1214_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1214",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1214_ack_0,
          idata => idata,
          odata => indvar350_1214,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1214
    phi_stmt_1408: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1411_wire & type_cast_1414_wire_constant;
      req <= phi_stmt_1408_req_0 & phi_stmt_1408_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1408",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1408_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1408,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1408
    phi_stmt_1453: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1457_wire_constant & type_cast_1459_wire;
      req <= phi_stmt_1453_req_0 & phi_stmt_1453_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1453",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1453_ack_0,
          idata => idata,
          odata => nx_x022x_xi295_1453,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1453
    phi_stmt_1460: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1464_wire_constant & type_cast_1466_wire;
      req <= phi_stmt_1460_req_0 & phi_stmt_1460_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1460",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1460_ack_0,
          idata => idata,
          odata => elementx_x021x_xi296_1460,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1460
    phi_stmt_1514: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1517_wire;
      req(0) <= phi_stmt_1514_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1514",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1514_ack_0,
          idata => idata,
          odata => shl8x_xi300x_xlcssa_1514,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1514
    phi_stmt_1624: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1627_wire & type_cast_1630_wire_constant;
      req <= phi_stmt_1624_req_0 & phi_stmt_1624_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1624",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1624_ack_0,
          idata => idata,
          odata => indvar_1624,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1624
    phi_stmt_745: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_749_wire_constant & type_cast_751_wire;
      req <= phi_stmt_745_req_0 & phi_stmt_745_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_745",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_745_ack_0,
          idata => idata,
          odata => indvar364_745,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_745
    phi_stmt_939: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_942_wire & type_cast_945_wire_constant;
      req <= phi_stmt_939_req_0 & phi_stmt_939_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_939",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_939_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_939,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_939
    phi_stmt_980: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_984_wire_constant & type_cast_986_wire;
      req <= phi_stmt_980_req_0 & phi_stmt_980_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_980",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_980_ack_0,
          idata => idata,
          odata => nx_x022x_xi_980,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_980
    phi_stmt_987: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_991_wire_constant & type_cast_993_wire;
      req <= phi_stmt_987_req_0 & phi_stmt_987_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_987",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_987_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_987,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_987
    -- flow-through select operator MUX_1210_inst
    umax23_1211 <= tmp21_1198 when (tmp22_1204(0) /=  '0') else type_cast_1209_wire_constant;
    -- flow-through select operator MUX_1389_inst
    umax_1390 <= tmp345_1146 when (tmp346_1152(0) /=  '0') else type_cast_1388_wire_constant;
    -- flow-through select operator MUX_741_inst
    umax31_742 <= tmp29_729 when (tmp30_735(0) /=  '0') else type_cast_740_wire_constant;
    -- flow-through select operator MUX_920_inst
    umax360_921 <= tmp358_694 when (tmp359_700(0) /=  '0') else type_cast_919_wire_constant;
    addr_of_1074_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1074_final_reg_req_0;
      addr_of_1074_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1074_final_reg_req_1;
      addr_of_1074_final_reg_ack_1<= rack(0);
      addr_of_1074_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1074_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1073_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1075,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1227_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1227_final_reg_req_0;
      addr_of_1227_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1227_final_reg_req_1;
      addr_of_1227_final_reg_ack_1<= rack(0);
      addr_of_1227_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1227_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1226_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1547_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1547_final_reg_req_0;
      addr_of_1547_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1547_final_reg_req_1;
      addr_of_1547_final_reg_ack_1<= rack(0);
      addr_of_1547_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1547_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1546_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_1548,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_758_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_758_final_reg_req_0;
      addr_of_758_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_758_final_reg_req_1;
      addr_of_758_final_reg_ack_1<= rack(0);
      addr_of_758_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_758_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_757_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1012_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1012_inst_req_0;
      type_cast_1012_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1012_inst_req_1;
      type_cast_1012_inst_ack_1<= rack(0);
      type_cast_1012_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1012_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1009,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1013,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1027_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1027_inst_req_0;
      type_cast_1027_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1027_inst_req_1;
      type_cast_1027_inst_ack_1<= rack(0);
      type_cast_1027_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1027_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1000,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1028,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1044_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1044_inst_req_0;
      type_cast_1044_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1044_inst_req_1;
      type_cast_1044_inst_ack_1<= rack(0);
      type_cast_1044_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1044_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1024,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1044_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1084_inst_req_0;
      type_cast_1084_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1084_inst_req_1;
      type_cast_1084_inst_ack_1<= rack(0);
      type_cast_1084_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1084_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1085,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1088_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1088_inst_req_0;
      type_cast_1088_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1088_inst_req_1;
      type_cast_1088_inst_ack_1<= rack(0);
      type_cast_1088_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1088_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1089,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1092_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1092_inst_req_0;
      type_cast_1092_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1092_inst_req_1;
      type_cast_1092_inst_ack_1<= rack(0);
      type_cast_1092_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1092_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_1093,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1096_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1096_inst_req_0;
      type_cast_1096_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1096_inst_req_1;
      type_cast_1096_inst_ack_1<= rack(0);
      type_cast_1096_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1096_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1097,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1121_inst
    process(sext_1118) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1118(63 downto 0);
      type_cast_1121_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1126_inst
    process(ASHR_i64_i64_1125_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1125_wire(63 downto 0);
      conv155_1127 <= tmp_var; -- 
    end process;
    type_cast_1155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1155_inst_req_0;
      type_cast_1155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1155_inst_req_1;
      type_cast_1155_inst_ack_1<= rack(0);
      type_cast_1155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_1156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1159_inst_req_0;
      type_cast_1159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1159_inst_req_1;
      type_cast_1159_inst_ack_1<= rack(0);
      type_cast_1159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1168_inst_req_0;
      type_cast_1168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1168_inst_req_1;
      type_cast_1168_inst_ack_1<= rack(0);
      type_cast_1168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1177_inst_req_0;
      type_cast_1177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1177_inst_req_1;
      type_cast_1177_inst_ack_1<= rack(0);
      type_cast_1177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp17_1178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1186_inst_req_0;
      type_cast_1186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1186_inst_req_1;
      type_cast_1186_inst_ack_1<= rack(0);
      type_cast_1186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp18_1183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_1187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1191_inst_req_0;
      type_cast_1191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1191_inst_req_1;
      type_cast_1191_inst_ack_1<= rack(0);
      type_cast_1191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1190_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1192,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1220_inst_req_0;
      type_cast_1220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1220_inst_req_1;
      type_cast_1220_inst_ack_1<= rack(0);
      type_cast_1220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext351_1371,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1220_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1234_inst_req_0;
      type_cast_1234_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1234_inst_req_1;
      type_cast_1234_inst_ack_1<= rack(0);
      type_cast_1234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1231,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1247_inst_req_0;
      type_cast_1247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1247_inst_req_1;
      type_cast_1247_inst_ack_1<= rack(0);
      type_cast_1247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1265_inst_req_0;
      type_cast_1265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1265_inst_req_1;
      type_cast_1265_inst_ack_1<= rack(0);
      type_cast_1265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1283_inst_req_0;
      type_cast_1283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1283_inst_req_1;
      type_cast_1283_inst_ack_1<= rack(0);
      type_cast_1283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1301_inst_req_0;
      type_cast_1301_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1301_inst_req_1;
      type_cast_1301_inst_ack_1<= rack(0);
      type_cast_1301_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1301_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1302,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1319_inst_req_0;
      type_cast_1319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1319_inst_req_1;
      type_cast_1319_inst_ack_1<= rack(0);
      type_cast_1319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1337_inst_req_0;
      type_cast_1337_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1337_inst_req_1;
      type_cast_1337_inst_ack_1<= rack(0);
      type_cast_1337_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1337_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_1334,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_1338,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1355_inst_req_0;
      type_cast_1355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1355_inst_req_1;
      type_cast_1355_inst_ack_1<= rack(0);
      type_cast_1355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_1352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_1356,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1399_inst
    process(tmp347_1396) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp347_1396(63 downto 0);
      type_cast_1399_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1404_inst
    process(ASHR_i64_i64_1403_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1403_wire(63 downto 0);
      phitmp325_1405 <= tmp_var; -- 
    end process;
    type_cast_1411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1411_inst_req_0;
      type_cast_1411_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1411_inst_req_1;
      type_cast_1411_inst_ack_1<= rack(0);
      type_cast_1411_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1411_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp325_1405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1411_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1443_inst_req_0;
      type_cast_1443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1443_inst_req_1;
      type_cast_1443_inst_ack_1<= rack(0);
      type_cast_1443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_54_1440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi292_1444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1459_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1459_inst_req_0;
      type_cast_1459_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1459_inst_req_1;
      type_cast_1459_inst_ack_1<= rack(0);
      type_cast_1459_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1459_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_62_1479,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1459_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1466_inst_req_0;
      type_cast_1466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1466_inst_req_1;
      type_cast_1466_inst_ack_1<= rack(0);
      type_cast_1466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi300_1497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1466_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1485_inst_req_0;
      type_cast_1485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1485_inst_req_1;
      type_cast_1485_inst_ack_1<= rack(0);
      type_cast_1485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi297_1482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi298_1486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1500_inst_req_0;
      type_cast_1500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1500_inst_req_1;
      type_cast_1500_inst_ack_1<= rack(0);
      type_cast_1500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp326_1473,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi301_1501,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1517_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1517_inst_req_0;
      type_cast_1517_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1517_inst_req_1;
      type_cast_1517_inst_ack_1<= rack(0);
      type_cast_1517_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1517_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi300_1497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1517_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1596_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1596_inst_req_0;
      type_cast_1596_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1596_inst_req_1;
      type_cast_1596_inst_ack_1<= rack(0);
      type_cast_1596_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1596_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp327_1593,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1597,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1606_inst_req_0;
      type_cast_1606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1606_inst_req_1;
      type_cast_1606_inst_ack_1<= rack(0);
      type_cast_1606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1615_inst_req_0;
      type_cast_1615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1615_inst_req_1;
      type_cast_1615_inst_ack_1<= rack(0);
      type_cast_1615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_1612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1627_inst_req_0;
      type_cast_1627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1627_inst_req_1;
      type_cast_1627_inst_ack_1<= rack(0);
      type_cast_1627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1627_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1644_inst_req_0;
      type_cast_1644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1644_inst_req_1;
      type_cast_1644_inst_ack_1<= rack(0);
      type_cast_1644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul254_1636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1648_inst_req_0;
      type_cast_1648_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1648_inst_req_1;
      type_cast_1648_inst_ack_1<= rack(0);
      type_cast_1648_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1648_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul260_1641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv261_1649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1681_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1681_inst_req_0;
      type_cast_1681_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1681_inst_req_1;
      type_cast_1681_inst_ack_1<= rack(0);
      type_cast_1681_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1681_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1680_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_1682,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1689_inst_req_0;
      type_cast_1689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1689_inst_req_1;
      type_cast_1689_inst_ack_1<= rack(0);
      type_cast_1689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1688_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv285_1690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_442_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_442_inst_req_0;
      type_cast_442_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_442_inst_req_1;
      type_cast_442_inst_ack_1<= rack(0);
      type_cast_442_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_442_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_439,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_443,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_455_inst_req_0;
      type_cast_455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_455_inst_req_1;
      type_cast_455_inst_ack_1<= rack(0);
      type_cast_455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_467_inst_req_0;
      type_cast_467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_467_inst_req_1;
      type_cast_467_inst_ack_1<= rack(0);
      type_cast_467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_468,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_480_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_480_inst_req_0;
      type_cast_480_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_480_inst_req_1;
      type_cast_480_inst_ack_1<= rack(0);
      type_cast_480_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_480_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_477,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_481,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_492_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_492_inst_req_0;
      type_cast_492_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_492_inst_req_1;
      type_cast_492_inst_ack_1<= rack(0);
      type_cast_492_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_492_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_505_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_505_inst_req_0;
      type_cast_505_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_505_inst_req_1;
      type_cast_505_inst_ack_1<= rack(0);
      type_cast_505_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_505_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_502,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_506,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_517_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_517_inst_req_0;
      type_cast_517_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_517_inst_req_1;
      type_cast_517_inst_ack_1<= rack(0);
      type_cast_517_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_517_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_514,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_518,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_530_inst_req_0;
      type_cast_530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_530_inst_req_1;
      type_cast_530_inst_ack_1<= rack(0);
      type_cast_530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_530_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_527,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_531,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_542_inst_req_0;
      type_cast_542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_542_inst_req_1;
      type_cast_542_inst_ack_1<= rack(0);
      type_cast_542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_542_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_555_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_555_inst_req_0;
      type_cast_555_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_555_inst_req_1;
      type_cast_555_inst_ack_1<= rack(0);
      type_cast_555_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_555_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_552,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_556,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_567_inst_req_0;
      type_cast_567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_567_inst_req_1;
      type_cast_567_inst_ack_1<= rack(0);
      type_cast_567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_564,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_568,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_580_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_580_inst_req_0;
      type_cast_580_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_580_inst_req_1;
      type_cast_580_inst_ack_1<= rack(0);
      type_cast_580_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_580_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_581,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_592_inst_req_1;
      type_cast_592_inst_ack_1<= rack(0);
      type_cast_592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_605_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_605_inst_req_0;
      type_cast_605_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_605_inst_req_1;
      type_cast_605_inst_ack_1<= rack(0);
      type_cast_605_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_605_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_606,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_617_inst_req_0;
      type_cast_617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_617_inst_req_1;
      type_cast_617_inst_ack_1<= rack(0);
      type_cast_617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_617_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_630_inst_req_0;
      type_cast_630_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_630_inst_req_1;
      type_cast_630_inst_ack_1<= rack(0);
      type_cast_630_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_630_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_639_inst_req_0;
      type_cast_639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_639_inst_req_1;
      type_cast_639_inst_ack_1<= rack(0);
      type_cast_639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_486,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_643_inst_req_0;
      type_cast_643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_643_inst_req_1;
      type_cast_643_inst_ack_1<= rack(0);
      type_cast_643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_659_inst_req_0;
      type_cast_659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_659_inst_req_1;
      type_cast_659_inst_ack_1<= rack(0);
      type_cast_659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_658_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_660,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_687_inst_req_0;
      type_cast_687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_687_inst_req_1;
      type_cast_687_inst_ack_1<= rack(0);
      type_cast_687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_686_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp357_688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_703_inst_req_0;
      type_cast_703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_703_inst_req_1;
      type_cast_703_inst_ack_1<= rack(0);
      type_cast_703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_703_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_486,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_704,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_712_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_712_inst_req_0;
      type_cast_712_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_712_inst_req_1;
      type_cast_712_inst_ack_1<= rack(0);
      type_cast_712_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_712_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp26_713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_722_inst_req_0;
      type_cast_722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_722_inst_req_1;
      type_cast_722_inst_ack_1<= rack(0);
      type_cast_722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_721_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp28_723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_751_inst_req_1;
      type_cast_751_inst_ack_1<= rack(0);
      type_cast_751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext365_902,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_751_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_765_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_765_inst_req_0;
      type_cast_765_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_765_inst_req_1;
      type_cast_765_inst_ack_1<= rack(0);
      type_cast_765_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_765_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_762,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_766,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_778_inst_req_0;
      type_cast_778_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_778_inst_req_1;
      type_cast_778_inst_ack_1<= rack(0);
      type_cast_778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_775,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_796_inst_req_0;
      type_cast_796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_796_inst_req_1;
      type_cast_796_inst_ack_1<= rack(0);
      type_cast_796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_796_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_814_inst_req_0;
      type_cast_814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_814_inst_req_1;
      type_cast_814_inst_ack_1<= rack(0);
      type_cast_814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_814_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_832_inst_req_0;
      type_cast_832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_832_inst_req_1;
      type_cast_832_inst_ack_1<= rack(0);
      type_cast_832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_850_inst_req_0;
      type_cast_850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_850_inst_req_1;
      type_cast_850_inst_ack_1<= rack(0);
      type_cast_850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_868_inst_req_0;
      type_cast_868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_868_inst_req_1;
      type_cast_868_inst_ack_1<= rack(0);
      type_cast_868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_865,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_869,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_886_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_886_inst_req_0;
      type_cast_886_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_886_inst_req_1;
      type_cast_886_inst_ack_1<= rack(0);
      type_cast_886_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_886_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_883,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_887,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_930_inst
    process(tmp361_927) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp361_927(63 downto 0);
      type_cast_930_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_935_inst
    process(ASHR_i64_i64_934_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_934_wire(63 downto 0);
      phitmp_936 <= tmp_var; -- 
    end process;
    type_cast_942_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_942_inst_req_0;
      type_cast_942_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_942_inst_req_1;
      type_cast_942_inst_ack_1<= rack(0);
      type_cast_942_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_942_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_936,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_942_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_986_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_986_inst_req_0;
      type_cast_986_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_986_inst_req_1;
      type_cast_986_inst_ack_1<= rack(0);
      type_cast_986_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_986_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_34_1006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_986_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_993_inst_req_0;
      type_cast_993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_993_inst_req_1;
      type_cast_993_inst_ack_1<= rack(0);
      type_cast_993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1024,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1073_index_1_rename
    process(R_ix_x0x_xlcssa_1072_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1072_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1072_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1073_index_1_resize
    process(ix_x0x_xlcssa_939) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_939;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1072_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1073_root_address_inst
    process(array_obj_ref_1073_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1073_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1073_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1226_index_1_rename
    process(R_indvar350_1225_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar350_1225_resized;
      ov(13 downto 0) := iv;
      R_indvar350_1225_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1226_index_1_resize
    process(indvar350_1214) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar350_1214;
      ov := iv(13 downto 0);
      R_indvar350_1225_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1226_root_address_inst
    process(array_obj_ref_1226_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1226_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1226_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1546_index_1_rename
    process(R_ix_x1x_xlcssa_1545_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1545_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1545_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1546_index_1_resize
    process(ix_x1x_xlcssa_1408) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1408;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1545_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1546_root_address_inst
    process(array_obj_ref_1546_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1546_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1546_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_757_index_1_rename
    process(R_indvar364_756_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar364_756_resized;
      ov(13 downto 0) := iv;
      R_indvar364_756_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_757_index_1_resize
    process(indvar364_745) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar364_745;
      ov := iv(13 downto 0);
      R_indvar364_756_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_757_root_address_inst
    process(array_obj_ref_757_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_757_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_757_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1077_addr_0
    process(ptr_deref_1077_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1077_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1077_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1077_base_resize
    process(arrayidx143_1075) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1075;
      ov := iv(13 downto 0);
      ptr_deref_1077_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1077_gather_scatter
    process(shl14x_xi_1068) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1068;
      ov(63 downto 0) := iv;
      ptr_deref_1077_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1077_root_address_inst
    process(ptr_deref_1077_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1077_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1077_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1363_addr_0
    process(ptr_deref_1363_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1363_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1363_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1363_base_resize
    process(arrayidx211_1228) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1228;
      ov := iv(13 downto 0);
      ptr_deref_1363_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1363_gather_scatter
    process(add207_1361) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_1361;
      ov(63 downto 0) := iv;
      ptr_deref_1363_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1363_root_address_inst
    process(ptr_deref_1363_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1363_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1363_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1550_addr_0
    process(ptr_deref_1550_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1550_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1550_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1550_base_resize
    process(arrayidx226_1548) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_1548;
      ov := iv(13 downto 0);
      ptr_deref_1550_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1550_gather_scatter
    process(shl14x_xi310_1541) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi310_1541;
      ov(63 downto 0) := iv;
      ptr_deref_1550_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1550_root_address_inst
    process(ptr_deref_1550_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1550_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1550_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_894_addr_0
    process(ptr_deref_894_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_894_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_894_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_894_base_resize
    process(arrayidx_759) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_759;
      ov := iv(13 downto 0);
      ptr_deref_894_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_894_gather_scatter
    process(add132_892) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_892;
      ov(63 downto 0) := iv;
      ptr_deref_894_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_894_root_address_inst
    process(ptr_deref_894_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_894_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_894_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1034_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1033;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1034_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1034_branch_req_0,
          ack0 => if_stmt_1034_branch_ack_0,
          ack1 => if_stmt_1034_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1134_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161317_1133;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1134_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1134_branch_req_0,
          ack0 => if_stmt_1134_branch_ack_0,
          ack1 => if_stmt_1134_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1377_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1376;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1377_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1377_branch_req_0,
          ack0 => if_stmt_1377_branch_ack_0,
          ack1 => if_stmt_1377_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1428_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_1427;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1428_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1428_branch_req_0,
          ack0 => if_stmt_1428_branch_ack_0,
          ack1 => if_stmt_1428_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1507_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi302_1506;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1507_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1507_branch_req_0,
          ack0 => if_stmt_1507_branch_ack_0,
          ack1 => if_stmt_1507_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1671_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1670;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1671_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1671_branch_req_0,
          ack0 => if_stmt_1671_branch_ack_0,
          ack1 => if_stmt_1671_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_667_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp321_666;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_667_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_667_branch_req_0,
          ack0 => if_stmt_667_branch_ack_0,
          ack1 => if_stmt_667_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_908_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond32_907;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_908_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_908_branch_req_0,
          ack0 => if_stmt_908_branch_ack_0,
          ack1 => if_stmt_908_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_959_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_958;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_959_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_959_branch_req_0,
          ack0 => if_stmt_959_branch_ack_0,
          ack1 => if_stmt_959_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1005_inst
    process(nx_x022x_xi_980) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_980, type_cast_1004_wire_constant, tmp_var);
      iNsTr_34_1006 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1472_inst
    process(nx_x022x_xi295_1453) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi295_1453, type_cast_1471_wire_constant, tmp_var);
      tmp326_1473 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1478_inst
    process(nx_x022x_xi295_1453) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi295_1453, type_cast_1477_wire_constant, tmp_var);
      iNsTr_62_1479 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1580_inst
    process(add43_561) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43_561, type_cast_1579_wire_constant, tmp_var);
      sub_1581 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1586_inst
    process(add63_611) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add63_611, type_cast_1585_wire_constant, tmp_var);
      sub269_1587 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1592_inst
    process(add53_586) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_586, type_cast_1591_wire_constant, tmp_var);
      tmp327_1593 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_999_inst
    process(nx_x022x_xi_980) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_980, type_cast_998_wire_constant, tmp_var);
      tmp_1000 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1602_inst
    process(tmp3_1597) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1597, type_cast_1601_wire_constant, tmp_var);
      tmp4_1603 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1640_inst
    process(tmp9_1621, mul254_1636) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_1621, mul254_1636, tmp_var);
      mul260_1641 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1664_inst
    process(indvar_1624) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1624, type_cast_1663_wire_constant, tmp_var);
      indvarx_xnext_1665 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1370_inst
    process(indvar350_1214) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar350_1214, type_cast_1369_wire_constant, tmp_var);
      indvarx_xnext351_1371 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_901_inst
    process(indvar364_745) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar364_745, type_cast_900_wire_constant, tmp_var);
      indvarx_xnext365_902 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1449_inst
    process(conv2x_xi292_1444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi292_1444, type_cast_1448_wire_constant, tmp_var);
      shlx_xi293_1450 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_976_inst
    process(conv2x_xi_971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_971, type_cast_975_wire_constant, tmp_var);
      shlx_xi_977 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1056_inst
    process(Bx_xnot_1051) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1051, type_cast_1055_wire_constant, tmp_var);
      add1216x_xi_1057 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1420_inst
    process(conv155_1127) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1127, type_cast_1419_wire_constant, tmp_var);
      and217_1421 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1529_inst
    process(iNsTr_70_1524) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_70_1524, type_cast_1528_wire_constant, tmp_var);
      add1216x_xi308_1530 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_951_inst
    process(conv83_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_660, type_cast_950_wire_constant, tmp_var);
      and_952 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1125_inst
    process(type_cast_1121_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1121_wire, type_cast_1124_wire_constant, tmp_var);
      ASHR_i64_i64_1125_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1403_inst
    process(type_cast_1399_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1399_wire, type_cast_1402_wire_constant, tmp_var);
      ASHR_i64_i64_1403_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_934_inst
    process(type_cast_930_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_930_wire, type_cast_933_wire_constant, tmp_var);
      ASHR_i64_i64_934_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1669_inst
    process(indvarx_xnext_1665, tmp4_1603) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1665, tmp4_1603, tmp_var);
      exitcond5_1670 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1375_inst
    process(indvarx_xnext351_1371, umax23_1211) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext351_1371, umax23_1211, tmp_var);
      exitcond_1376 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1426_inst
    process(and217_1421) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_1421, type_cast_1425_wire_constant, tmp_var);
      tobool218_1427 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_906_inst
    process(indvarx_xnext365_902, umax31_742) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext365_902, umax31_742, tmp_var);
      exitcond32_907 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_957_inst
    process(and_952) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_952, type_cast_956_wire_constant, tmp_var);
      tobool_958 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1145_inst
    process(conv155_1127) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1127, type_cast_1144_wire_constant, tmp_var);
      tmp345_1146 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1197_inst
    process(tmp20_1192) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1192, type_cast_1196_wire_constant, tmp_var);
      tmp21_1198 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_693_inst
    process(tmp357_688) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp357_688, type_cast_692_wire_constant, tmp_var);
      tmp358_694 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_728_inst
    process(tmp28_723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp28_723, type_cast_727_wire_constant, tmp_var);
      tmp29_729 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1562_inst
    process(add73_636, add23_511) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_636, add23_511, tmp_var);
      mul236_1563 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1567_inst
    process(add43_561, add33_536) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add43_561, add33_536, tmp_var);
      mul249_1568 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1611_inst
    process(add73_636, add23_511) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_636, add23_511, tmp_var);
      tmp7_1612 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1620_inst
    process(tmp6_1607, tmp8_1616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_1607, tmp8_1616, tmp_var);
      tmp9_1621 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1635_inst
    process(tmp9_1621, indvar_1624) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1621, indvar_1624, tmp_var);
      mul254_1636 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_648_inst
    process(conv79_640, add_461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_640, add_461, tmp_var);
      mul_649 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_653_inst
    process(mul_649, conv81_644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_649, conv81_644, tmp_var);
      mul82_654 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_677_inst
    process(add_461, conv79_640) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_461, conv79_640, tmp_var);
      tmp354_678 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_682_inst
    process(tmp354_678, conv81_644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp354_678, conv81_644, tmp_var);
      tmp356_683 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_708_inst
    process(add_461, tmp24_704) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_461, tmp24_704, tmp_var);
      tmp25_709 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_717_inst
    process(tmp25_709, tmp26_713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_709, tmp26_713, tmp_var);
      tmp27_718 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1101_inst
    process(conv153_1097, conv145_1085) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1097, conv145_1085, tmp_var);
      mul148_1102 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1106_inst
    process(mul148_1102, conv150_1093) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1102, conv150_1093, tmp_var);
      mul151_1107 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1111_inst
    process(mul151_1107, conv147_1089) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1107, conv147_1089, tmp_var);
      mul154_1112 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1164_inst
    process(tmp12_1156, tmp13_1160) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1156, tmp13_1160, tmp_var);
      tmp14_1165 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1173_inst
    process(tmp14_1165, tmp15_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1165, tmp15_1169, tmp_var);
      tmp16_1174 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1182_inst
    process(tmp16_1174, tmp17_1178) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_1174, tmp17_1178, tmp_var);
      tmp18_1183 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_485_inst
    process(shl10_474, conv12_481) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_474, conv12_481, tmp_var);
      add13_486 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_510_inst
    process(shl20_499, conv22_506) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_499, conv22_506, tmp_var);
      add23_511 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_535_inst
    process(shl30_524, conv32_531) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_524, conv32_531, tmp_var);
      add33_536 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_560_inst
    process(shl40_549, conv42_556) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_549, conv42_556, tmp_var);
      add43_561 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_585_inst
    process(shl50_574, conv52_581) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_574, conv52_581, tmp_var);
      add53_586 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_610_inst
    process(shl60_599, conv62_606) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_599, conv62_606, tmp_var);
      add63_611 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_635_inst
    process(shl70_624, conv72_631) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_624, conv72_631, tmp_var);
      add73_636 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_460_inst
    process(shl_449, conv3_456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_449, conv3_456, tmp_var);
      add_461 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1017_inst
    process(conv5x_xi_1013, elementx_x021x_xi_987) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1013, elementx_x021x_xi_987, tmp_var);
      addx_xi_1018 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1252_inst
    process(shl167_1241, conv170_1248) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1241, conv170_1248, tmp_var);
      add171_1253 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1270_inst
    process(shl173_1259, conv176_1266) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1259, conv176_1266, tmp_var);
      add177_1271 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1288_inst
    process(shl179_1277, conv182_1284) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1277, conv182_1284, tmp_var);
      add183_1289 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1306_inst
    process(shl185_1295, conv188_1302) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1295, conv188_1302, tmp_var);
      add189_1307 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1324_inst
    process(shl191_1313, conv194_1320) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1313, conv194_1320, tmp_var);
      add195_1325 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1342_inst
    process(shl197_1331, conv200_1338) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_1331, conv200_1338, tmp_var);
      add201_1343 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1360_inst
    process(shl203_1349, conv206_1356) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_1349, conv206_1356, tmp_var);
      add207_1361 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1490_inst
    process(conv5x_xi298_1486, elementx_x021x_xi296_1460) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi298_1486, elementx_x021x_xi296_1460, tmp_var);
      addx_xi299_1491 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_783_inst
    process(shl92_772, conv95_779) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_772, conv95_779, tmp_var);
      add96_784 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_801_inst
    process(shl98_790, conv101_797) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_790, conv101_797, tmp_var);
      add102_802 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_819_inst
    process(shl104_808, conv107_815) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_808, conv107_815, tmp_var);
      add108_820 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_837_inst
    process(shl110_826, conv113_833) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_826, conv113_833, tmp_var);
      add114_838 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_855_inst
    process(shl116_844, conv119_851) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_844, conv119_851, tmp_var);
      add120_856 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_873_inst
    process(shl122_862, conv125_869) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_862, conv125_869, tmp_var);
      add126_874 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_891_inst
    process(shl128_880, conv131_887) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_880, conv131_887, tmp_var);
      add132_892 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_473_inst
    process(conv9_468) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_468, type_cast_472_wire_constant, tmp_var);
      shl10_474 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_498_inst
    process(conv19_493) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_493, type_cast_497_wire_constant, tmp_var);
      shl20_499 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_523_inst
    process(conv29_518) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_518, type_cast_522_wire_constant, tmp_var);
      shl30_524 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_548_inst
    process(conv39_543) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_543, type_cast_547_wire_constant, tmp_var);
      shl40_549 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_573_inst
    process(conv49_568) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_568, type_cast_572_wire_constant, tmp_var);
      shl50_574 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_598_inst
    process(conv59_593) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_593, type_cast_597_wire_constant, tmp_var);
      shl60_599 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_623_inst
    process(conv69_618) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_618, type_cast_622_wire_constant, tmp_var);
      shl70_624 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_448_inst
    process(conv1_443) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_443, type_cast_447_wire_constant, tmp_var);
      shl_449 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_970_inst
    process(mul82_654) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_654, type_cast_969_wire_constant, tmp_var);
      conv2x_xi_971 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1023_inst
    process(addx_xi_1018) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1018, type_cast_1022_wire_constant, tmp_var);
      shl8x_xi_1024 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1050_inst
    process(conv83_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_660, type_cast_1049_wire_constant, tmp_var);
      Bx_xnot_1051 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1067_inst
    process(shl8x_xix_xlcssa_1041, sh_promx_xi_1063) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1041, sh_promx_xi_1063, tmp_var);
      shl14x_xi_1068 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1117_inst
    process(mul154_1112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1112, type_cast_1116_wire_constant, tmp_var);
      sext_1118 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1240_inst
    process(conv165_1235) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1235, type_cast_1239_wire_constant, tmp_var);
      shl167_1241 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1258_inst
    process(add171_1253) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1253, type_cast_1257_wire_constant, tmp_var);
      shl173_1259 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1276_inst
    process(add177_1271) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1271, type_cast_1275_wire_constant, tmp_var);
      shl179_1277 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1294_inst
    process(add183_1289) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1289, type_cast_1293_wire_constant, tmp_var);
      shl185_1295 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1312_inst
    process(add189_1307) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1307, type_cast_1311_wire_constant, tmp_var);
      shl191_1313 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1330_inst
    process(add195_1325) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_1325, type_cast_1329_wire_constant, tmp_var);
      shl197_1331 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1348_inst
    process(add201_1343) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_1343, type_cast_1347_wire_constant, tmp_var);
      shl203_1349 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1395_inst
    process(umax_1390) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1390, type_cast_1394_wire_constant, tmp_var);
      tmp347_1396 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1439_inst
    process(mul154_1112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1112, type_cast_1438_wire_constant, tmp_var);
      iNsTr_54_1440 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1496_inst
    process(addx_xi299_1491) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi299_1491, type_cast_1495_wire_constant, tmp_var);
      shl8x_xi300_1497 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1523_inst
    process(mul154_1112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1112, type_cast_1522_wire_constant, tmp_var);
      iNsTr_70_1524 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1540_inst
    process(shl8x_xi300x_xlcssa_1514, sh_promx_xi309_1536) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi300x_xlcssa_1514, sh_promx_xi309_1536, tmp_var);
      shl14x_xi310_1541 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_771_inst
    process(conv90_766) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_766, type_cast_770_wire_constant, tmp_var);
      shl92_772 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_789_inst
    process(add96_784) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_784, type_cast_788_wire_constant, tmp_var);
      shl98_790 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_807_inst
    process(add102_802) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_802, type_cast_806_wire_constant, tmp_var);
      shl104_808 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_825_inst
    process(add108_820) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_820, type_cast_824_wire_constant, tmp_var);
      shl110_826 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_843_inst
    process(add114_838) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_838, type_cast_842_wire_constant, tmp_var);
      shl116_844 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_861_inst
    process(add120_856) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_856, type_cast_860_wire_constant, tmp_var);
      shl122_862 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_879_inst
    process(add126_874) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_874, type_cast_878_wire_constant, tmp_var);
      shl128_880 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_926_inst
    process(umax360_921) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax360_921, type_cast_925_wire_constant, tmp_var);
      tmp361_927 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1694_inst
    process(conv285_1690, conv230_1682) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv285_1690, conv230_1682, tmp_var);
      sub289_1695 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_665_inst
    process(mul82_654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_654, type_cast_664_wire_constant, tmp_var);
      cmp321_666 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1132_inst
    process(conv155_1127) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1127, type_cast_1131_wire_constant, tmp_var);
      cmp161317_1133 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1151_inst
    process(tmp345_1146) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp345_1146, type_cast_1150_wire_constant, tmp_var);
      tmp346_1152 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1203_inst
    process(tmp21_1198) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp21_1198, type_cast_1202_wire_constant, tmp_var);
      tmp22_1204 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_699_inst
    process(tmp358_694) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp358_694, type_cast_698_wire_constant, tmp_var);
      tmp359_700 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_734_inst
    process(tmp29_729) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp29_729, type_cast_733_wire_constant, tmp_var);
      tmp30_735 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1032_inst
    process(convx_xi_1028, shlx_xi_977) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1028, shlx_xi_977, tmp_var);
      cmpx_xi_1033 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1505_inst
    process(convx_xi301_1501, shlx_xi293_1450) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi301_1501, shlx_xi293_1450, tmp_var);
      cmpx_xi302_1506 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1062_inst
    process(add1216x_xi_1057) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1057, type_cast_1061_wire_constant, tmp_var);
      sh_promx_xi_1063 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1535_inst
    process(add1216x_xi308_1530) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi308_1530, type_cast_1534_wire_constant, tmp_var);
      sh_promx_xi309_1536 <= tmp_var; --
    end process;
    -- shared split operator group (115) : array_obj_ref_1073_index_offset 
    ApIntAdd_group_115: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1072_scaled;
      array_obj_ref_1073_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1073_index_offset_req_0;
      array_obj_ref_1073_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1073_index_offset_req_1;
      array_obj_ref_1073_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_115_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_115_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_115",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 115
    -- shared split operator group (116) : array_obj_ref_1226_index_offset 
    ApIntAdd_group_116: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar350_1225_scaled;
      array_obj_ref_1226_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1226_index_offset_req_0;
      array_obj_ref_1226_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1226_index_offset_req_1;
      array_obj_ref_1226_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_116_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_116_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_116",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 116
    -- shared split operator group (117) : array_obj_ref_1546_index_offset 
    ApIntAdd_group_117: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1545_scaled;
      array_obj_ref_1546_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1546_index_offset_req_0;
      array_obj_ref_1546_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1546_index_offset_req_1;
      array_obj_ref_1546_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_117_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : array_obj_ref_757_index_offset 
    ApIntAdd_group_118: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar364_756_scaled;
      array_obj_ref_757_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_757_index_offset_req_0;
      array_obj_ref_757_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_757_index_offset_req_1;
      array_obj_ref_757_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_118_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- unary operator type_cast_1190_inst
    process(tmp19_1187) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp19_1187, tmp_var);
      type_cast_1190_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1680_inst
    process(call229_1557) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_1557, tmp_var);
      type_cast_1680_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1688_inst
    process(call284_1685) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call284_1685, tmp_var);
      type_cast_1688_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_658_inst
    process(mul82_654) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_654, tmp_var);
      type_cast_658_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_686_inst
    process(tmp356_683) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp356_683, tmp_var);
      type_cast_686_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_721_inst
    process(tmp27_718) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp27_718, tmp_var);
      type_cast_721_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_894_store_0 ptr_deref_1077_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_894_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1077_store_0_req_0;
      ptr_deref_894_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1077_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_894_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1077_store_0_req_1;
      ptr_deref_894_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1077_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_894_word_address_0 & ptr_deref_1077_word_address_0;
      data_in <= ptr_deref_894_data_0 & ptr_deref_1077_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1363_store_0 ptr_deref_1550_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1363_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1550_store_0_req_0;
      ptr_deref_1363_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1550_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1363_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1550_store_0_req_1;
      ptr_deref_1363_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1550_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1363_word_address_0 & ptr_deref_1550_word_address_0;
      data_in <= ptr_deref_1363_data_0 & ptr_deref_1550_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_761_inst RPIPE_maxpool_input_pipe_774_inst RPIPE_maxpool_input_pipe_792_inst RPIPE_maxpool_input_pipe_810_inst RPIPE_maxpool_input_pipe_828_inst RPIPE_maxpool_input_pipe_438_inst RPIPE_maxpool_input_pipe_451_inst RPIPE_maxpool_input_pipe_463_inst RPIPE_maxpool_input_pipe_476_inst RPIPE_maxpool_input_pipe_488_inst RPIPE_maxpool_input_pipe_501_inst RPIPE_maxpool_input_pipe_513_inst RPIPE_maxpool_input_pipe_526_inst RPIPE_maxpool_input_pipe_538_inst RPIPE_maxpool_input_pipe_551_inst RPIPE_maxpool_input_pipe_563_inst RPIPE_maxpool_input_pipe_576_inst RPIPE_maxpool_input_pipe_588_inst RPIPE_maxpool_input_pipe_601_inst RPIPE_maxpool_input_pipe_613_inst RPIPE_maxpool_input_pipe_626_inst RPIPE_maxpool_input_pipe_846_inst RPIPE_maxpool_input_pipe_864_inst RPIPE_maxpool_input_pipe_882_inst RPIPE_maxpool_input_pipe_1008_inst RPIPE_maxpool_input_pipe_1230_inst RPIPE_maxpool_input_pipe_1243_inst RPIPE_maxpool_input_pipe_1261_inst RPIPE_maxpool_input_pipe_1279_inst RPIPE_maxpool_input_pipe_1297_inst RPIPE_maxpool_input_pipe_1315_inst RPIPE_maxpool_input_pipe_1333_inst RPIPE_maxpool_input_pipe_1351_inst RPIPE_maxpool_input_pipe_1481_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_761_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_774_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_792_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_810_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_828_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_438_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_451_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_463_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_476_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_488_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_501_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_513_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_526_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_538_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_551_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_563_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_576_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_588_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_601_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_613_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_626_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_846_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_864_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_882_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1008_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1230_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1243_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1261_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1279_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1297_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1315_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1333_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1351_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1481_inst_req_0;
      RPIPE_maxpool_input_pipe_761_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_774_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_792_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_810_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_828_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_438_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_451_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_463_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_476_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_488_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_501_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_513_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_526_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_538_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_551_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_563_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_576_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_588_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_601_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_613_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_626_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_846_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_864_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_882_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1008_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1230_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1243_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1261_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1279_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1297_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1315_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1333_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1351_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1481_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_761_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_774_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_792_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_810_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_828_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_438_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_451_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_463_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_476_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_488_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_501_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_513_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_526_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_538_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_551_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_563_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_576_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_588_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_601_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_613_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_626_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_846_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_864_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_882_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1008_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1230_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1243_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1261_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1279_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1297_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1315_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1333_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1351_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1481_inst_req_1;
      RPIPE_maxpool_input_pipe_761_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_774_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_792_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_810_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_828_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_438_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_451_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_463_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_476_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_488_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_501_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_513_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_526_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_538_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_551_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_563_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_576_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_588_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_601_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_613_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_626_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_846_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_864_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_882_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1008_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1230_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1243_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1261_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1279_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1297_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1315_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1333_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1351_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1481_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call89_762 <= data_out(271 downto 264);
      call93_775 <= data_out(263 downto 256);
      call99_793 <= data_out(255 downto 248);
      call105_811 <= data_out(247 downto 240);
      call111_829 <= data_out(239 downto 232);
      call_439 <= data_out(231 downto 224);
      call2_452 <= data_out(223 downto 216);
      call6_464 <= data_out(215 downto 208);
      call11_477 <= data_out(207 downto 200);
      call16_489 <= data_out(199 downto 192);
      call21_502 <= data_out(191 downto 184);
      call26_514 <= data_out(183 downto 176);
      call31_527 <= data_out(175 downto 168);
      call36_539 <= data_out(167 downto 160);
      call41_552 <= data_out(159 downto 152);
      call46_564 <= data_out(151 downto 144);
      call51_577 <= data_out(143 downto 136);
      call56_589 <= data_out(135 downto 128);
      call61_602 <= data_out(127 downto 120);
      call66_614 <= data_out(119 downto 112);
      call71_627 <= data_out(111 downto 104);
      call117_847 <= data_out(103 downto 96);
      call123_865 <= data_out(95 downto 88);
      call129_883 <= data_out(87 downto 80);
      callx_xi_1009 <= data_out(79 downto 72);
      call164_1231 <= data_out(71 downto 64);
      call168_1244 <= data_out(63 downto 56);
      call174_1262 <= data_out(55 downto 48);
      call180_1280 <= data_out(47 downto 40);
      call186_1298 <= data_out(39 downto 32);
      call192_1316 <= data_out(31 downto 24);
      call198_1334 <= data_out(23 downto 16);
      call204_1352 <= data_out(15 downto 8);
      callx_xi297_1482 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1696_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1696_inst_req_0;
      WPIPE_elapsed_time_pipe_1696_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1696_inst_req_1;
      WPIPE_elapsed_time_pipe_1696_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub289_1695;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_1572_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1572_inst_req_0;
      WPIPE_maxpool_output_pipe_1572_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1572_inst_req_1;
      WPIPE_maxpool_output_pipe_1572_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1574_wire_constant;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_num_out_pipe_1569_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1569_inst_req_0;
      WPIPE_num_out_pipe_1569_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1569_inst_req_1;
      WPIPE_num_out_pipe_1569_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul249_1568;
      num_out_pipe_write_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_1557_call call_stmt_1685_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1557_call_req_0;
      reqL_unguarded(0) <= call_stmt_1685_call_req_0;
      call_stmt_1557_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1685_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1557_call_req_1;
      reqR_unguarded(0) <= call_stmt_1685_call_req_1;
      call_stmt_1557_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1685_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_1557 <= data_out(127 downto 64);
      call284_1685 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1652_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1652_call_req_0;
      call_stmt_1652_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1652_call_req_1;
      call_stmt_1652_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv255_1645 & conv261_1649;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(127 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1659_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1659_call_req_0;
      call_stmt_1659_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1659_call_req_1;
      call_stmt_1659_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul236_1563 & add33_536 & sub_1581 & sub269_1587 & add23_511 & add13_486;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_3814_start: Boolean;
  signal convolve_CP_3814_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nacc_1778_1730_buf_req_0 : boolean;
  signal nacc_1778_1730_buf_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1745_inst_ack_0 : boolean;
  signal n_out_count_1807_1735_buf_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1745_inst_ack_1 : boolean;
  signal nacc_1778_1730_buf_req_1 : boolean;
  signal nacc_1778_1730_buf_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_1745_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1745_inst_req_0 : boolean;
  signal phi_stmt_1731_ack_0 : boolean;
  signal phi_stmt_1731_req_0 : boolean;
  signal n_out_count_1807_1735_buf_req_0 : boolean;
  signal n_out_count_1807_1735_buf_ack_0 : boolean;
  signal n_out_count_1807_1735_buf_ack_1 : boolean;
  signal phi_stmt_1731_req_1 : boolean;
  signal RPIPE_input_pipe1_1738_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1738_inst_ack_1 : boolean;
  signal RPIPE_input_pipe1_1738_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1738_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1707_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1707_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1707_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1707_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1710_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1710_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1710_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1710_inst_ack_1 : boolean;
  signal do_while_stmt_1721_branch_req_0 : boolean;
  signal phi_stmt_1723_req_1 : boolean;
  signal phi_stmt_1723_req_0 : boolean;
  signal phi_stmt_1723_ack_0 : boolean;
  signal nmycount_1786_1726_buf_req_0 : boolean;
  signal nmycount_1786_1726_buf_ack_0 : boolean;
  signal nmycount_1786_1726_buf_req_1 : boolean;
  signal nmycount_1786_1726_buf_ack_1 : boolean;
  signal phi_stmt_1727_req_1 : boolean;
  signal phi_stmt_1727_req_0 : boolean;
  signal phi_stmt_1727_ack_0 : boolean;
  signal SUB_u32_u32_1759_inst_req_0 : boolean;
  signal SUB_u32_u32_1759_inst_ack_0 : boolean;
  signal SUB_u32_u32_1759_inst_req_1 : boolean;
  signal SUB_u32_u32_1759_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_1793_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1793_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1793_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_1793_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1814_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_1814_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_1814_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1814_inst_ack_1 : boolean;
  signal slice_1819_inst_req_0 : boolean;
  signal slice_1819_inst_ack_0 : boolean;
  signal slice_1819_inst_req_1 : boolean;
  signal slice_1819_inst_ack_1 : boolean;
  signal slice_1823_inst_req_0 : boolean;
  signal slice_1823_inst_ack_0 : boolean;
  signal slice_1823_inst_req_1 : boolean;
  signal slice_1823_inst_ack_1 : boolean;
  signal W_next_sum_1801_delayed_1_0_1825_inst_req_0 : boolean;
  signal W_next_sum_1801_delayed_1_0_1825_inst_ack_0 : boolean;
  signal W_next_sum_1801_delayed_1_0_1825_inst_req_1 : boolean;
  signal W_next_sum_1801_delayed_1_0_1825_inst_ack_1 : boolean;
  signal type_cast_1831_inst_req_0 : boolean;
  signal type_cast_1831_inst_ack_0 : boolean;
  signal type_cast_1831_inst_req_1 : boolean;
  signal type_cast_1831_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1829_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1829_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1829_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1829_inst_ack_1 : boolean;
  signal W_next_sum_1806_delayed_1_0_1833_inst_req_0 : boolean;
  signal W_next_sum_1806_delayed_1_0_1833_inst_ack_0 : boolean;
  signal W_next_sum_1806_delayed_1_0_1833_inst_req_1 : boolean;
  signal W_next_sum_1806_delayed_1_0_1833_inst_ack_1 : boolean;
  signal type_cast_1839_inst_req_0 : boolean;
  signal type_cast_1839_inst_ack_0 : boolean;
  signal type_cast_1839_inst_req_1 : boolean;
  signal type_cast_1839_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_ack_1 : boolean;
  signal do_while_stmt_1721_branch_ack_0 : boolean;
  signal do_while_stmt_1721_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_3814_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3814_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_3814_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3814_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_3814: Block -- control-path 
    signal convolve_CP_3814_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convolve_CP_3814_elements(0) <= convolve_CP_3814_start;
    convolve_CP_3814_symbol <= convolve_CP_3814_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1705/$entry
      -- CP-element group 0: 	 branch_block_stmt_1705/branch_block_stmt_1705__entry__
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720__entry__
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/$entry
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Sample/rr
      -- 
    rr_3836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(0), ack => RPIPE_num_out_pipe_1707_inst_req_0); -- 
    rr_3850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(0), ack => RPIPE_size_pipe_1710_inst_req_0); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1705/$exit
      -- CP-element group 1: 	 branch_block_stmt_1705/branch_block_stmt_1705__exit__
      -- CP-element group 1: 	 branch_block_stmt_1705/do_while_stmt_1721__exit__
      -- 
    convolve_CP_3814_elements(1) <= convolve_CP_3814_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Update/cr
      -- 
    ra_3837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1707_inst_ack_0, ack => convolve_CP_3814_elements(2)); -- 
    cr_3841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(2), ack => RPIPE_num_out_pipe_1707_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_num_out_pipe_1707_Update/ca
      -- 
    ca_3842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1707_inst_ack_1, ack => convolve_CP_3814_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Update/cr
      -- 
    ra_3851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1710_inst_ack_0, ack => convolve_CP_3814_elements(4)); -- 
    cr_3855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(4), ack => RPIPE_size_pipe_1710_inst_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/RPIPE_size_pipe_1710_Update/ca
      -- 
    ca_3856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1710_inst_ack_1, ack => convolve_CP_3814_elements(5)); -- 
    -- CP-element group 6:  join  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720__exit__
      -- CP-element group 6: 	 branch_block_stmt_1705/do_while_stmt_1721__entry__
      -- CP-element group 6: 	 branch_block_stmt_1705/assign_stmt_1708_to_assign_stmt_1720/$exit
      -- 
    convolve_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "convolve_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(3) & convolve_CP_3814_elements(5);
      gj_convolve_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1705/do_while_stmt_1721/$entry
      -- CP-element group 7: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721__entry__
      -- 
    convolve_CP_3814_elements(7) <= convolve_CP_3814_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	127 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721__exit__
      -- 
    -- Element group convolve_CP_3814_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_back
      -- 
    -- Element group convolve_CP_3814_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	125 
    -- CP-element group 10: 	126 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1705/do_while_stmt_1721/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_taken/$entry
      -- 
    convolve_CP_3814_elements(10) <= convolve_CP_3814_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	124 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_body_done
      -- 
    convolve_CP_3814_elements(11) <= convolve_CP_3814_elements(124);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	24 
    -- CP-element group 12: 	43 
    -- CP-element group 12: 	62 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_3814_elements(12) <= convolve_CP_3814_elements(9);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	45 
    -- CP-element group 13: 	64 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_3814_elements(13) <= convolve_CP_3814_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	83 
    -- CP-element group 14: 	123 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_3814_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	123 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/condition_evaluated
      -- 
    condition_evaluated_3871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(15), ack => do_while_stmt_1721_branch_req_0); -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(19) & convolve_CP_3814_elements(123);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	37 
    -- CP-element group 16: 	56 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	58 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_sample_start__ps
      -- 
    convolve_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(20) & convolve_CP_3814_elements(37) & convolve_CP_3814_elements(56) & convolve_CP_3814_elements(19);
      gj_convolve_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	59 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	76 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	84 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	37 
    -- CP-element group 17: 	56 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_sample_completed_
      -- 
    convolve_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(22) & convolve_CP_3814_elements(40) & convolve_CP_3814_elements(59);
      gj_convolve_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	57 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	60 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_update_start__ps
      -- 
    convolve_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(21) & convolve_CP_3814_elements(38) & convolve_CP_3814_elements(57);
      gj_convolve_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	61 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(23) & convolve_CP_3814_elements(42) & convolve_CP_3814_elements(61);
      gj_convolve_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	86 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_sample_start_
      -- 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(17) & convolve_CP_3814_elements(86);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	103 
    -- CP-element group 21: 	114 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_update_start_
      -- 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(91) & convolve_CP_3814_elements(103) & convolve_CP_3814_elements(114);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_sample_completed__ps
      -- 
    -- Element group convolve_CP_3814_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: 	90 
    -- CP-element group 23: 	101 
    -- CP-element group 23: 	112 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_update_completed__ps
      -- 
    -- Element group convolve_CP_3814_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	12 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_loopback_trigger
      -- 
    convolve_CP_3814_elements(24) <= convolve_CP_3814_elements(12);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_loopback_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_loopback_sample_req_ps
      -- 
    phi_stmt_1723_loopback_sample_req_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1723_loopback_sample_req_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(25), ack => phi_stmt_1723_req_1); -- 
    -- Element group convolve_CP_3814_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_entry_trigger
      -- 
    convolve_CP_3814_elements(26) <= convolve_CP_3814_elements(13);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_entry_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_entry_sample_req_ps
      -- 
    phi_stmt_1723_entry_sample_req_3889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1723_entry_sample_req_3889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(27), ack => phi_stmt_1723_req_0); -- 
    -- Element group convolve_CP_3814_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_phi_mux_ack
      -- CP-element group 28: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1723_phi_mux_ack_ps
      -- 
    phi_stmt_1723_phi_mux_ack_3892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1723_ack_0, ack => convolve_CP_3814_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_sample_completed_
      -- 
    -- Element group convolve_CP_3814_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_update_start_
      -- 
    -- Element group convolve_CP_3814_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_update_completed__ps
      -- 
    convolve_CP_3814_elements(31) <= convolve_CP_3814_elements(32);
    -- CP-element group 32:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	31 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_mcount_var_1725_update_completed_
      -- 
    -- Element group convolve_CP_3814_elements(32) is a control-delay.
    cp_element_32_delay: control_delay_element  generic map(name => " 32_delay", delay_value => 1)  port map(req => convolve_CP_3814_elements(30), ack => convolve_CP_3814_elements(32), clk => clk, reset =>reset);
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Sample/req
      -- 
    req_3913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(33), ack => nmycount_1786_1726_buf_req_0); -- 
    -- Element group convolve_CP_3814_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Update/req
      -- 
    req_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(34), ack => nmycount_1786_1726_buf_req_1); -- 
    -- Element group convolve_CP_3814_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Sample/ack
      -- 
    ack_3914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1786_1726_buf_ack_0, ack => convolve_CP_3814_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nmycount_1726_Update/ack
      -- 
    ack_3919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1786_1726_buf_ack_1, ack => convolve_CP_3814_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	17 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	16 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_sample_start_
      -- 
    convolve_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(17) & convolve_CP_3814_elements(78) & convolve_CP_3814_elements(82) & convolve_CP_3814_elements(86);
      gj_convolve_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	95 
    -- CP-element group 38: 	99 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	18 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_update_start_
      -- 
    convolve_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(95) & convolve_CP_3814_elements(99);
      gj_convolve_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_sample_start__ps
      -- 
    convolve_CP_3814_elements(39) <= convolve_CP_3814_elements(16);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	17 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_sample_completed__ps
      -- 
    -- Element group convolve_CP_3814_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_update_start__ps
      -- 
    convolve_CP_3814_elements(41) <= convolve_CP_3814_elements(18);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: 	93 
    -- CP-element group 42: 	97 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_update_completed__ps
      -- 
    -- Element group convolve_CP_3814_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	12 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_loopback_trigger
      -- 
    convolve_CP_3814_elements(43) <= convolve_CP_3814_elements(12);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_loopback_sample_req_ps
      -- 
    phi_stmt_1727_loopback_sample_req_3930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1727_loopback_sample_req_3930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(44), ack => phi_stmt_1727_req_1); -- 
    -- Element group convolve_CP_3814_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	13 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_entry_trigger
      -- 
    convolve_CP_3814_elements(45) <= convolve_CP_3814_elements(13);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_entry_sample_req_ps
      -- 
    phi_stmt_1727_entry_sample_req_3933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1727_entry_sample_req_3933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(46), ack => phi_stmt_1727_req_0); -- 
    -- Element group convolve_CP_3814_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1727_phi_mux_ack_ps
      -- 
    phi_stmt_1727_phi_mux_ack_3936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1727_ack_0, ack => convolve_CP_3814_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_sample_start_
      -- 
    -- Element group convolve_CP_3814_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_update_start__ps
      -- 
    -- Element group convolve_CP_3814_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_update_completed__ps
      -- 
    convolve_CP_3814_elements(50) <= convolve_CP_3814_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_acc_var_1729_update_completed_
      -- 
    -- Element group convolve_CP_3814_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => convolve_CP_3814_elements(49), ack => convolve_CP_3814_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Sample/$entry
      -- 
    req_3957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(52), ack => nacc_1778_1730_buf_req_0); -- 
    -- Element group convolve_CP_3814_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Update/req
      -- CP-element group 53: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_update_start_
      -- 
    req_3962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(53), ack => nacc_1778_1730_buf_req_1); -- 
    -- Element group convolve_CP_3814_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Sample/$exit
      -- 
    ack_3958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1778_1730_buf_ack_0, ack => convolve_CP_3814_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_nacc_1730_update_completed__ps
      -- 
    ack_3963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1778_1730_buf_ack_1, ack => convolve_CP_3814_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	17 
    -- CP-element group 56: 	86 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	16 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_sample_start_
      -- 
    convolve_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(17) & convolve_CP_3814_elements(86);
      gj_convolve_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	88 
    -- CP-element group 57: 	91 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	18 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_update_start_
      -- 
    convolve_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(88) & convolve_CP_3814_elements(91);
      gj_convolve_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_sample_start__ps
      -- 
    convolve_CP_3814_elements(58) <= convolve_CP_3814_elements(16);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_sample_completed__ps
      -- 
    -- Element group convolve_CP_3814_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	18 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_update_start__ps
      -- 
    convolve_CP_3814_elements(60) <= convolve_CP_3814_elements(18);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	87 
    -- CP-element group 61: 	90 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_update_completed__ps
      -- 
    -- Element group convolve_CP_3814_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	12 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_loopback_trigger
      -- 
    convolve_CP_3814_elements(62) <= convolve_CP_3814_elements(12);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_loopback_sample_req_ps
      -- 
    phi_stmt_1731_loopback_sample_req_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1731_loopback_sample_req_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(63), ack => phi_stmt_1731_req_1); -- 
    -- Element group convolve_CP_3814_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	13 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_entry_trigger
      -- 
    convolve_CP_3814_elements(64) <= convolve_CP_3814_elements(13);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_entry_sample_req_ps
      -- CP-element group 65: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_entry_sample_req
      -- 
    phi_stmt_1731_entry_sample_req_3977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1731_entry_sample_req_3977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(65), ack => phi_stmt_1731_req_0); -- 
    -- Element group convolve_CP_3814_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_phi_mux_ack
      -- CP-element group 66: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/phi_stmt_1731_phi_mux_ack_ps
      -- 
    phi_stmt_1731_phi_mux_ack_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1731_ack_0, ack => convolve_CP_3814_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_sample_start_
      -- 
    -- Element group convolve_CP_3814_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_update_start_
      -- CP-element group 68: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_update_start__ps
      -- 
    -- Element group convolve_CP_3814_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_update_completed__ps
      -- 
    convolve_CP_3814_elements(69) <= convolve_CP_3814_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1734_update_completed_
      -- 
    -- Element group convolve_CP_3814_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convolve_CP_3814_elements(68), ack => convolve_CP_3814_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_sample_start__ps
      -- CP-element group 71: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Sample/$entry
      -- 
    req_4001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(71), ack => n_out_count_1807_1735_buf_req_0); -- 
    -- Element group convolve_CP_3814_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_update_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Update/req
      -- CP-element group 72: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Update/$entry
      -- 
    req_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(72), ack => n_out_count_1807_1735_buf_req_1); -- 
    -- Element group convolve_CP_3814_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_sample_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Sample/$exit
      -- 
    ack_4002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1807_1735_buf_ack_0, ack => convolve_CP_3814_elements(73)); -- 
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_update_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/R_n_out_count_1735_Update/$exit
      -- 
    ack_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1807_1735_buf_ack_1, ack => convolve_CP_3814_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	78 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Sample/rr
      -- 
    rr_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(75), ack => RPIPE_input_pipe1_1738_inst_req_0); -- 
    convolve_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(78);
      gj_convolve_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	17 
    -- CP-element group 76: 	77 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	95 
    -- CP-element group 76: 	99 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_update_start_
      -- CP-element group 76: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Update/cr
      -- 
    cr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(76), ack => RPIPE_input_pipe1_1738_inst_req_1); -- 
    convolve_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(17) & convolve_CP_3814_elements(77) & convolve_CP_3814_elements(95) & convolve_CP_3814_elements(99);
      gj_convolve_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	76 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Sample/ra
      -- 
    ra_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1738_inst_ack_0, ack => convolve_CP_3814_elements(77)); -- 
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	97 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	75 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_input_pipe1_1738_update_completed_
      -- 
    ca_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1738_inst_ack_1, ack => convolve_CP_3814_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Sample/$entry
      -- 
    rr_4030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(79), ack => RPIPE_kernel_pipe1_1745_inst_req_0); -- 
    convolve_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(82);
      gj_convolve_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: 	81 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	88 
    -- CP-element group 80: 	95 
    -- CP-element group 80: 	99 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_update_start_
      -- CP-element group 80: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Update/$entry
      -- 
    cr_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(80), ack => RPIPE_kernel_pipe1_1745_inst_req_1); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(17) & convolve_CP_3814_elements(81) & convolve_CP_3814_elements(88) & convolve_CP_3814_elements(95) & convolve_CP_3814_elements(99);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Sample/$exit
      -- 
    ra_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1745_inst_ack_0, ack => convolve_CP_3814_elements(81)); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	87 
    -- CP-element group 82: 	93 
    -- CP-element group 82: 	97 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/RPIPE_kernel_pipe1_1745_Update/ca
      -- 
    ca_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1745_inst_ack_1, ack => convolve_CP_3814_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	14 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Sample/rr
      -- 
    rr_4044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(83), ack => SUB_u32_u32_1759_inst_req_0); -- 
    convolve_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(14) & convolve_CP_3814_elements(85);
      gj_convolve_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	17 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	91 
    -- CP-element group 84: 	103 
    -- CP-element group 84: 	114 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Update/cr
      -- 
    cr_4049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(84), ack => SUB_u32_u32_1759_inst_req_1); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(17) & convolve_CP_3814_elements(91) & convolve_CP_3814_elements(103) & convolve_CP_3814_elements(114);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Sample/ra
      -- 
    ra_4045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1759_inst_ack_0, ack => convolve_CP_3814_elements(85)); -- 
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	90 
    -- CP-element group 86: 	101 
    -- CP-element group 86: 	112 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	20 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	56 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/SUB_u32_u32_1759_Update/ca
      -- 
    ca_4050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1759_inst_ack_1, ack => convolve_CP_3814_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	61 
    -- CP-element group 87: 	82 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Sample/req
      -- 
    req_4058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(87), ack => WPIPE_kernel_pipe1_1793_inst_req_0); -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(61) & convolve_CP_3814_elements(82) & convolve_CP_3814_elements(89);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	57 
    -- CP-element group 88: 	80 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Sample/ack
      -- CP-element group 88: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Update/req
      -- 
    ack_4059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1793_inst_ack_0, ack => convolve_CP_3814_elements(88)); -- 
    req_4063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(88), ack => WPIPE_kernel_pipe1_1793_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	124 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_kernel_pipe1_1793_Update/ack
      -- 
    ack_4064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1793_inst_ack_1, ack => convolve_CP_3814_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	23 
    -- CP-element group 90: 	61 
    -- CP-element group 90: 	86 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Sample/req
      -- 
    req_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(90), ack => WPIPE_input_done_pipe_1814_inst_req_0); -- 
    convolve_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(23) & convolve_CP_3814_elements(61) & convolve_CP_3814_elements(86) & convolve_CP_3814_elements(92);
      gj_convolve_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	21 
    -- CP-element group 91: 	57 
    -- CP-element group 91: 	84 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Update/req
      -- 
    ack_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1814_inst_ack_0, ack => convolve_CP_3814_elements(91)); -- 
    req_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(91), ack => WPIPE_input_done_pipe_1814_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	124 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_input_done_pipe_1814_Update/ack
      -- 
    ack_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1814_inst_ack_1, ack => convolve_CP_3814_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	42 
    -- CP-element group 93: 	78 
    -- CP-element group 93: 	82 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Sample/rr
      -- 
    rr_4086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(93), ack => slice_1819_inst_req_0); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(42) & convolve_CP_3814_elements(78) & convolve_CP_3814_elements(82) & convolve_CP_3814_elements(95);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	107 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Update/cr
      -- 
    cr_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(94), ack => slice_1819_inst_req_1); -- 
    convolve_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3814_elements(107);
      gj_convolve_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	38 
    -- CP-element group 95: 	76 
    -- CP-element group 95: 	80 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Sample/ra
      -- 
    ra_4087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1819_inst_ack_0, ack => convolve_CP_3814_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1819_Update/ca
      -- 
    ca_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1819_inst_ack_1, ack => convolve_CP_3814_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	42 
    -- CP-element group 97: 	78 
    -- CP-element group 97: 	82 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Sample/rr
      -- 
    rr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(97), ack => slice_1823_inst_req_0); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(42) & convolve_CP_3814_elements(78) & convolve_CP_3814_elements(82) & convolve_CP_3814_elements(99);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	118 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Update/cr
      -- 
    cr_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(98), ack => slice_1823_inst_req_1); -- 
    convolve_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3814_elements(118);
      gj_convolve_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	38 
    -- CP-element group 99: 	76 
    -- CP-element group 99: 	80 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Sample/ra
      -- 
    ra_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1823_inst_ack_0, ack => convolve_CP_3814_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	116 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/slice_1823_Update/ca
      -- 
    ca_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1823_inst_ack_1, ack => convolve_CP_3814_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	23 
    -- CP-element group 101: 	86 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Sample/req
      -- 
    req_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(101), ack => W_next_sum_1801_delayed_1_0_1825_inst_req_0); -- 
    convolve_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(23) & convolve_CP_3814_elements(86) & convolve_CP_3814_elements(103);
      gj_convolve_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: 	110 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Update/req
      -- 
    req_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(102), ack => W_next_sum_1801_delayed_1_0_1825_inst_req_1); -- 
    convolve_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(107) & convolve_CP_3814_elements(110);
      gj_convolve_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	21 
    -- CP-element group 103: 	84 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Sample/ack
      -- 
    ack_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1801_delayed_1_0_1825_inst_ack_0, ack => convolve_CP_3814_elements(103)); -- 
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	109 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1827_Update/ack
      -- 
    ack_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1801_delayed_1_0_1825_inst_ack_1, ack => convolve_CP_3814_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	96 
    -- CP-element group 105: 	104 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Sample/rr
      -- 
    rr_4128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(105), ack => type_cast_1831_inst_req_0); -- 
    convolve_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(96) & convolve_CP_3814_elements(104) & convolve_CP_3814_elements(107);
      gj_convolve_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	110 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_update_start_
      -- CP-element group 106: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Update/cr
      -- 
    cr_4133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(106), ack => type_cast_1831_inst_req_1); -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3814_elements(110);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	94 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Sample/ra
      -- 
    ra_4129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_0, ack => convolve_CP_3814_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1831_Update/ca
      -- 
    ca_4134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_1, ack => convolve_CP_3814_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	104 
    -- CP-element group 109: 	108 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	122 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Sample/req
      -- 
    req_4142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(109), ack => WPIPE_maxpool_output_pipe_1829_inst_req_0); -- 
    convolve_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(104) & convolve_CP_3814_elements(108) & convolve_CP_3814_elements(122);
      gj_convolve_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	102 
    -- CP-element group 110: 	106 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Sample/ack
      -- CP-element group 110: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Update/req
      -- 
    ack_4143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1829_inst_ack_0, ack => convolve_CP_3814_elements(110)); -- 
    req_4147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(110), ack => WPIPE_maxpool_output_pipe_1829_inst_req_1); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	120 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1829_Update/ack
      -- 
    ack_4148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1829_inst_ack_1, ack => convolve_CP_3814_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	23 
    -- CP-element group 112: 	86 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Sample/req
      -- 
    req_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(112), ack => W_next_sum_1806_delayed_1_0_1833_inst_req_0); -- 
    convolve_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(23) & convolve_CP_3814_elements(86) & convolve_CP_3814_elements(114);
      gj_convolve_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	118 
    -- CP-element group 113: 	121 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Update/req
      -- 
    req_4161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(113), ack => W_next_sum_1806_delayed_1_0_1833_inst_req_1); -- 
    convolve_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(118) & convolve_CP_3814_elements(121);
      gj_convolve_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	21 
    -- CP-element group 114: 	84 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Sample/ack
      -- 
    ack_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1806_delayed_1_0_1833_inst_ack_0, ack => convolve_CP_3814_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/assign_stmt_1835_Update/ack
      -- 
    ack_4162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1806_delayed_1_0_1833_inst_ack_1, ack => convolve_CP_3814_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	100 
    -- CP-element group 116: 	115 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Sample/rr
      -- 
    rr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(116), ack => type_cast_1839_inst_req_0); -- 
    convolve_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(100) & convolve_CP_3814_elements(115) & convolve_CP_3814_elements(118);
      gj_convolve_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_update_start_
      -- CP-element group 117: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Update/cr
      -- 
    cr_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(117), ack => type_cast_1839_inst_req_1); -- 
    convolve_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3814_elements(121);
      gj_convolve_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	98 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Sample/ra
      -- 
    ra_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1839_inst_ack_0, ack => convolve_CP_3814_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/type_cast_1839_Update/ca
      -- 
    ca_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1839_inst_ack_1, ack => convolve_CP_3814_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	119 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Sample/req
      -- 
    req_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(120), ack => WPIPE_maxpool_output_pipe_1837_inst_req_0); -- 
    convolve_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(111) & convolve_CP_3814_elements(115) & convolve_CP_3814_elements(119) & convolve_CP_3814_elements(122);
      gj_convolve_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	113 
    -- CP-element group 121: 	117 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_update_start_
      -- CP-element group 121: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Sample/ack
      -- CP-element group 121: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Update/req
      -- 
    ack_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1837_inst_ack_0, ack => convolve_CP_3814_elements(121)); -- 
    req_4189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3814_elements(121), ack => WPIPE_maxpool_output_pipe_1837_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	109 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/WPIPE_maxpool_output_pipe_1837_Update/ack
      -- 
    ack_4190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1837_inst_ack_1, ack => convolve_CP_3814_elements(122)); -- 
    -- CP-element group 123:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	14 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	15 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_3814_elements(123) is a control-delay.
    cp_element_123_delay: control_delay_element  generic map(name => " 123_delay", delay_value => 1)  port map(req => convolve_CP_3814_elements(14), ack => convolve_CP_3814_elements(123), clk => clk, reset =>reset);
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	89 
    -- CP-element group 124: 	92 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	11 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1705/do_while_stmt_1721/do_while_stmt_1721_loop_body/$exit
      -- 
    convolve_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3814_elements(89) & convolve_CP_3814_elements(92) & convolve_CP_3814_elements(122);
      gj_convolve_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3814_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	10 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_exit/$exit
      -- CP-element group 125: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_exit/ack
      -- 
    ack_4195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1721_branch_ack_0, ack => convolve_CP_3814_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	10 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_taken/$exit
      -- CP-element group 126: 	 branch_block_stmt_1705/do_while_stmt_1721/loop_taken/ack
      -- 
    ack_4199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1721_branch_ack_1, ack => convolve_CP_3814_elements(126)); -- 
    -- CP-element group 127:  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	8 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1705/do_while_stmt_1721/$exit
      -- 
    convolve_CP_3814_elements(127) <= convolve_CP_3814_elements(8);
    convolve_do_while_stmt_1721_terminator_4200: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1721_terminator_4200", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_3814_elements(11),loop_continue => convolve_CP_3814_elements(126),loop_terminate => convolve_CP_3814_elements(125),loop_back => convolve_CP_3814_elements(9),loop_exit => convolve_CP_3814_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1723_phi_seq_3920_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3814_elements(26);
      convolve_CP_3814_elements(29)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3814_elements(29);
      convolve_CP_3814_elements(30)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3814_elements(31);
      convolve_CP_3814_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3814_elements(24);
      convolve_CP_3814_elements(33)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3814_elements(35);
      convolve_CP_3814_elements(34)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3814_elements(36);
      convolve_CP_3814_elements(25) <= phi_mux_reqs(1);
      phi_stmt_1723_phi_seq_3920 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1723_phi_seq_3920") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3814_elements(16), 
          phi_sample_ack => convolve_CP_3814_elements(22), 
          phi_update_req => convolve_CP_3814_elements(18), 
          phi_update_ack => convolve_CP_3814_elements(23), 
          phi_mux_ack => convolve_CP_3814_elements(28), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1727_phi_seq_3964_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3814_elements(45);
      convolve_CP_3814_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3814_elements(48);
      convolve_CP_3814_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3814_elements(50);
      convolve_CP_3814_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3814_elements(43);
      convolve_CP_3814_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3814_elements(54);
      convolve_CP_3814_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3814_elements(55);
      convolve_CP_3814_elements(44) <= phi_mux_reqs(1);
      phi_stmt_1727_phi_seq_3964 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1727_phi_seq_3964") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3814_elements(39), 
          phi_sample_ack => convolve_CP_3814_elements(40), 
          phi_update_req => convolve_CP_3814_elements(41), 
          phi_update_ack => convolve_CP_3814_elements(42), 
          phi_mux_ack => convolve_CP_3814_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1731_phi_seq_4008_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3814_elements(64);
      convolve_CP_3814_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3814_elements(67);
      convolve_CP_3814_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3814_elements(69);
      convolve_CP_3814_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3814_elements(62);
      convolve_CP_3814_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3814_elements(73);
      convolve_CP_3814_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3814_elements(74);
      convolve_CP_3814_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1731_phi_seq_4008 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1731_phi_seq_4008") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3814_elements(58), 
          phi_sample_ack => convolve_CP_3814_elements(59), 
          phi_update_req => convolve_CP_3814_elements(60), 
          phi_update_ack => convolve_CP_3814_elements(61), 
          phi_mux_ack => convolve_CP_3814_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3872_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_3814_elements(12);
        preds(1)  <= convolve_CP_3814_elements(13);
        entry_tmerge_3872 : transition_merge -- 
          generic map(name => " entry_tmerge_3872")
          port map (preds => preds, symbol_out => convolve_CP_3814_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1803_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_1784_wire : std_logic_vector(31 downto 0);
    signal MUX_1804_wire : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_1739_1739_delayed_1_0_1760 : std_logic_vector(31 downto 0);
    signal acc_1727 : std_logic_vector(15 downto 0);
    signal acc_val_1772 : std_logic_vector(15 downto 0);
    signal acc_val_dn_1824 : std_logic_vector(7 downto 0);
    signal acc_val_up_1820 : std_logic_vector(7 downto 0);
    signal acc_var_1720 : std_logic_vector(15 downto 0);
    signal all_done_flag_1812 : std_logic_vector(0 downto 0);
    signal iread_1739 : std_logic_vector(15 downto 0);
    signal ival_1743 : std_logic_vector(15 downto 0);
    signal konst_1758_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1775_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1781_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1783_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1802_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1815_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1842_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1746 : std_logic_vector(15 downto 0);
    signal kval_1750 : std_logic_vector(15 downto 0);
    signal mcount_var_1715 : std_logic_vector(31 downto 0);
    signal mul_val_1755 : std_logic_vector(15 downto 0);
    signal mycount_1723 : std_logic_vector(31 downto 0);
    signal n_out_count_1807 : std_logic_vector(15 downto 0);
    signal n_out_count_1807_1735_buffered : std_logic_vector(15 downto 0);
    signal nacc_1778 : std_logic_vector(15 downto 0);
    signal nacc_1778_1730_buffered : std_logic_vector(15 downto 0);
    signal next_sum_1765 : std_logic_vector(0 downto 0);
    signal next_sum_1801_delayed_1_0_1827 : std_logic_vector(0 downto 0);
    signal next_sum_1806_delayed_1_0_1835 : std_logic_vector(0 downto 0);
    signal nmycount_1786 : std_logic_vector(31 downto 0);
    signal nmycount_1786_1726_buffered : std_logic_vector(31 downto 0);
    signal num_out_1708 : std_logic_vector(15 downto 0);
    signal out_count_1731 : std_logic_vector(15 downto 0);
    signal out_done_flag_1791 : std_logic_vector(0 downto 0);
    signal size_1711 : std_logic_vector(31 downto 0);
    signal type_cast_1734_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1768_wire : std_logic_vector(15 downto 0);
    signal type_cast_1770_wire : std_logic_vector(15 downto 0);
    signal type_cast_1800_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1831_wire : std_logic_vector(7 downto 0);
    signal type_cast_1839_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    acc_var_1720 <= "0000000000000000";
    konst_1758_wire_constant <= "00000000000000000000000000000001";
    konst_1775_wire_constant <= "0000000000000000";
    konst_1781_wire_constant <= "00000000000000000000000000000000";
    konst_1783_wire_constant <= "00000000000000000000000000000001";
    konst_1802_wire_constant <= "0000000000000001";
    konst_1815_wire_constant <= "1";
    konst_1842_wire_constant <= "1";
    mcount_var_1715 <= "00000000000000000000000000000000";
    type_cast_1734_wire_constant <= "0000000000000001";
    type_cast_1800_wire_constant <= "0000000000000001";
    phi_stmt_1723: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= mcount_var_1715 & nmycount_1786_1726_buffered;
      req <= phi_stmt_1723_req_0 & phi_stmt_1723_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1723",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1723_ack_0,
          idata => idata,
          odata => mycount_1723,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1723
    phi_stmt_1727: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= acc_var_1720 & nacc_1778_1730_buffered;
      req <= phi_stmt_1727_req_0 & phi_stmt_1727_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1727",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1727_ack_0,
          idata => idata,
          odata => acc_1727,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1727
    phi_stmt_1731: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1734_wire_constant & n_out_count_1807_1735_buffered;
      req <= phi_stmt_1731_req_0 & phi_stmt_1731_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1731",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1731_ack_0,
          idata => idata,
          odata => out_count_1731,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1731
    -- flow-through select operator MUX_1777_inst
    nacc_1778 <= konst_1775_wire_constant when (next_sum_1765(0) /=  '0') else acc_val_1772;
    -- flow-through select operator MUX_1785_inst
    nmycount_1786 <= konst_1781_wire_constant when (next_sum_1765(0) /=  '0') else ADD_u32_u32_1784_wire;
    -- flow-through select operator MUX_1804_inst
    MUX_1804_wire <= type_cast_1800_wire_constant when (out_done_flag_1791(0) /=  '0') else ADD_u16_u16_1803_wire;
    -- flow-through select operator MUX_1806_inst
    n_out_count_1807 <= MUX_1804_wire when (next_sum_1765(0) /=  '0') else out_count_1731;
    slice_1819_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1819_inst_req_0;
      slice_1819_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1819_inst_req_1;
      slice_1819_inst_ack_1<= update_ack(0);
      slice_1819_inst: SliceSplitProtocol generic map(name => "slice_1819_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1772, dout => acc_val_up_1820, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1823_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1823_inst_req_0;
      slice_1823_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1823_inst_req_1;
      slice_1823_inst_ack_1<= update_ack(0);
      slice_1823_inst: SliceSplitProtocol generic map(name => "slice_1823_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1772, dout => acc_val_dn_1824, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_next_sum_1801_delayed_1_0_1825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1801_delayed_1_0_1825_inst_req_0;
      W_next_sum_1801_delayed_1_0_1825_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1801_delayed_1_0_1825_inst_req_1;
      W_next_sum_1801_delayed_1_0_1825_inst_ack_1<= rack(0);
      W_next_sum_1801_delayed_1_0_1825_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1801_delayed_1_0_1825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1801_delayed_1_0_1827,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_next_sum_1806_delayed_1_0_1833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1806_delayed_1_0_1833_inst_req_0;
      W_next_sum_1806_delayed_1_0_1833_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1806_delayed_1_0_1833_inst_req_1;
      W_next_sum_1806_delayed_1_0_1833_inst_ack_1<= rack(0);
      W_next_sum_1806_delayed_1_0_1833_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1806_delayed_1_0_1833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1806_delayed_1_0_1835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_out_count_1807_1735_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1807_1735_buf_req_0;
      n_out_count_1807_1735_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1807_1735_buf_req_1;
      n_out_count_1807_1735_buf_ack_1<= rack(0);
      n_out_count_1807_1735_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1807_1735_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1807_1735_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_1778_1730_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1778_1730_buf_req_0;
      nacc_1778_1730_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1778_1730_buf_req_1;
      nacc_1778_1730_buf_ack_1<= rack(0);
      nacc_1778_1730_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1778_1730_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1778_1730_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_1786_1726_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1786_1726_buf_req_0;
      nmycount_1786_1726_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1786_1726_buf_req_1;
      nmycount_1786_1726_buf_ack_1<= rack(0);
      nmycount_1786_1726_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1786_1726_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1786_1726_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1742_inst
    process(iread_1739) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1739(15 downto 0);
      ival_1743 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1749_inst
    process(kread_1746) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1746(15 downto 0);
      kval_1750 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1768_inst
    process(acc_1727) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := acc_1727(15 downto 0);
      type_cast_1768_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1770_inst
    process(mul_val_1755) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1755(15 downto 0);
      type_cast_1770_wire <= tmp_var; -- 
    end process;
    type_cast_1831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1831_inst_req_0;
      type_cast_1831_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1831_inst_req_1;
      type_cast_1831_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1801_delayed_1_0_1827(0);
      type_cast_1831_inst_gI: SplitGuardInterface generic map(name => "type_cast_1831_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_1820,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1831_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1839_inst_req_0;
      type_cast_1839_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1839_inst_req_1;
      type_cast_1839_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1806_delayed_1_0_1835(0);
      type_cast_1839_inst_gI: SplitGuardInterface generic map(name => "type_cast_1839_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_1824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1839_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1721_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1842_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1721_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1721_branch_req_0,
          ack0 => do_while_stmt_1721_branch_ack_0,
          ack1 => do_while_stmt_1721_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_1771_inst
    process(type_cast_1768_wire, type_cast_1770_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1768_wire, type_cast_1770_wire, tmp_var);
      acc_val_1772 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1803_inst
    process(out_count_1731) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1731, konst_1802_wire_constant, tmp_var);
      ADD_u16_u16_1803_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1784_inst
    process(mycount_1723) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1723, konst_1783_wire_constant, tmp_var);
      ADD_u32_u32_1784_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1811_inst
    process(out_done_flag_1791, next_sum_1765) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1791, next_sum_1765, tmp_var);
      all_done_flag_1812 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1790_inst
    process(out_count_1731, num_out_1708) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1731, num_out_1708, tmp_var);
      out_done_flag_1791 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1764_inst
    process(mycount_1723, SUB_u32_u32_1739_1739_delayed_1_0_1760) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1723, SUB_u32_u32_1739_1739_delayed_1_0_1760, tmp_var);
      next_sum_1765 <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_1754_inst
    process(kval_1750, ival_1743) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1750, ival_1743, tmp_var);
      mul_val_1755 <= tmp_var; --
    end process;
    -- shared split operator group (7) : SUB_u32_u32_1759_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1711;
      SUB_u32_u32_1739_1739_delayed_1_0_1760 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_1759_inst_req_0;
      SUB_u32_u32_1759_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_1759_inst_req_1;
      SUB_u32_u32_1759_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared inport operator group (0) : RPIPE_input_pipe1_1738_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1738_inst_req_0;
      RPIPE_input_pipe1_1738_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1738_inst_req_1;
      RPIPE_input_pipe1_1738_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1739 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1745_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1745_inst_req_0;
      RPIPE_kernel_pipe1_1745_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1745_inst_req_1;
      RPIPE_kernel_pipe1_1745_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      kread_1746 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_num_out_pipe_1707_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1707_inst_req_0;
      RPIPE_num_out_pipe_1707_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1707_inst_req_1;
      RPIPE_num_out_pipe_1707_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1708 <= data_out(15 downto 0);
      num_out_pipe_read_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_2: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_size_pipe_1710_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1710_inst_req_0;
      RPIPE_size_pipe_1710_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1710_inst_req_1;
      RPIPE_size_pipe_1710_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_1711 <= data_out(31 downto 0);
      size_pipe_read_3_gI: SplitGuardInterface generic map(name => "size_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_3: InputPortRevised -- 
        generic map ( name => "size_pipe_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1814_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1814_inst_req_0;
      WPIPE_input_done_pipe_1814_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1814_inst_req_1;
      WPIPE_input_done_pipe_1814_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1812(0);
      data_in <= konst_1815_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1793_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1793_inst_req_0;
      WPIPE_kernel_pipe1_1793_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1793_inst_req_1;
      WPIPE_kernel_pipe1_1793_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not out_done_flag_1791(0);
      data_in <= kread_1746;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_maxpool_output_pipe_1829_inst WPIPE_maxpool_output_pipe_1837_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1829_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1837_inst_req_0;
      WPIPE_maxpool_output_pipe_1829_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1837_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1829_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1837_inst_req_1;
      WPIPE_maxpool_output_pipe_1829_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1837_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1806_delayed_1_0_1835(0);
      guard_vector(1)  <= next_sum_1801_delayed_1_0_1827(0);
      data_in <= type_cast_1831_wire & type_cast_1839_wire;
      maxpool_output_pipe_write_2_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 128)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_676_start: Boolean;
  signal loadKernelChannel_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_fn_394_delayed_13_0_408_inst_ack_0 : boolean;
  signal array_obj_ref_397_index_offset_ack_0 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_1 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_428_inst_req_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_1 : boolean;
  signal my_fetch_339_359_buf_ack_1 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_1 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_ack_1 : boolean;
  signal array_obj_ref_397_index_offset_req_1 : boolean;
  signal array_obj_ref_397_index_offset_ack_1 : boolean;
  signal WPIPE_size_pipe_428_inst_req_0 : boolean;
  signal my_fetch_339_359_buf_req_0 : boolean;
  signal my_fetch_339_359_buf_req_1 : boolean;
  signal phi_stmt_356_req_0 : boolean;
  signal type_cast_432_inst_ack_1 : boolean;
  signal ptr_deref_406_load_0_req_0 : boolean;
  signal phi_stmt_356_req_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_1 : boolean;
  signal type_cast_432_inst_req_0 : boolean;
  signal addr_of_398_final_reg_req_0 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_1 : boolean;
  signal type_cast_432_inst_ack_0 : boolean;
  signal addr_of_398_final_reg_ack_0 : boolean;
  signal nfetch_val_419_358_buf_req_0 : boolean;
  signal addr_of_398_final_reg_req_1 : boolean;
  signal addr_of_398_final_reg_ack_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_0 : boolean;
  signal array_obj_ref_397_index_offset_req_0 : boolean;
  signal ptr_deref_406_load_0_ack_0 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_0 : boolean;
  signal nfetch_val_419_358_buf_ack_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_0 : boolean;
  signal phi_stmt_356_ack_0 : boolean;
  signal type_cast_432_inst_req_1 : boolean;
  signal do_while_stmt_350_branch_ack_1 : boolean;
  signal my_fetch_339_359_buf_ack_0 : boolean;
  signal nfetch_val_419_358_buf_req_1 : boolean;
  signal nfetch_val_419_358_buf_ack_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_0 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_1 : boolean;
  signal array_obj_ref_333_index_offset_req_0 : boolean;
  signal array_obj_ref_333_index_offset_ack_0 : boolean;
  signal array_obj_ref_333_index_offset_req_1 : boolean;
  signal array_obj_ref_333_index_offset_ack_1 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_1 : boolean;
  signal addr_of_334_final_reg_req_0 : boolean;
  signal addr_of_334_final_reg_ack_0 : boolean;
  signal addr_of_334_final_reg_req_1 : boolean;
  signal addr_of_334_final_reg_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_0 : boolean;
  signal do_while_stmt_350_branch_ack_0 : boolean;
  signal ptr_deref_406_load_0_ack_1 : boolean;
  signal ptr_deref_406_load_0_req_1 : boolean;
  signal ptr_deref_338_load_0_req_0 : boolean;
  signal ptr_deref_338_load_0_ack_0 : boolean;
  signal ptr_deref_338_load_0_req_1 : boolean;
  signal ptr_deref_338_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_1 : boolean;
  signal do_while_stmt_350_branch_req_0 : boolean;
  signal phi_stmt_352_req_0 : boolean;
  signal phi_stmt_352_req_1 : boolean;
  signal phi_stmt_352_ack_0 : boolean;
  signal nmycount_374_354_buf_req_0 : boolean;
  signal nmycount_374_354_buf_ack_0 : boolean;
  signal nmycount_374_354_buf_req_1 : boolean;
  signal nmycount_374_354_buf_ack_1 : boolean;
  signal start_add_355_buf_req_0 : boolean;
  signal start_add_355_buf_ack_0 : boolean;
  signal start_add_355_buf_req_1 : boolean;
  signal start_add_355_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 128) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(tag_length + 127 downto 128) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 127 downto 128);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_676: Block -- control-path 
    signal loadKernelChannel_CP_676_elements: BooleanArray(94 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_676_elements(0) <= loadKernelChannel_CP_676_start;
    loadKernelChannel_CP_676_symbol <= loadKernelChannel_CP_676_elements(94);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resized_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_computed_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/rr
      -- 
    req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => addr_of_334_final_reg_req_1); -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => RPIPE_input_done_pipe_347_inst_req_0); -- 
    cr_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => ptr_deref_338_load_0_req_1); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_0); -- 
    req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/ack
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_start_
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_offset_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/req
      -- 
    ack_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(2)); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(2), ack => addr_of_334_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_completed_
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$exit
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/ack
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_completed_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_start_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_resized
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/rr
      -- 
    ack_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(4)); -- 
    rr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(4), ack => ptr_deref_338_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_completed_
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/ra
      -- 
    ra_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_completed_
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_ack
      -- 
    ca_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_completed_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_start_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/ra
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$entry
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/cr
      -- 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_0, ack => loadKernelChannel_CP_676_elements(7)); -- 
    cr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(7), ack => RPIPE_input_done_pipe_347_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_completed_
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$exit
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/ca
      -- 
    ca_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_1, ack => loadKernelChannel_CP_676_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_328_to_assign_stmt_348/$exit
      -- CP-element group 9: 	 branch_block_stmt_349/$entry
      -- CP-element group 9: 	 branch_block_stmt_349/branch_block_stmt_349__entry__
      -- CP-element group 9: 	 branch_block_stmt_349/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(8) & loadKernelChannel_CP_676_elements(6) & loadKernelChannel_CP_676_elements(1);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	90 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	91 
    -- CP-element group 10: 	92 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_update_start_
      -- CP-element group 10: 	 assign_stmt_433/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_sample_start_
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/rr
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_349/$exit
      -- CP-element group 10: 	 branch_block_stmt_349/branch_block_stmt_349__exit__
      -- CP-element group 10: 	 branch_block_stmt_349/do_while_stmt_350__exit__
      -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_0); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_1); -- 
    loadKernelChannel_CP_676_elements(10) <= loadKernelChannel_CP_676_elements(90);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/$entry
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_CP_676_elements(11) <= loadKernelChannel_CP_676_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	90 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__exit__
      -- 
    -- Element group loadKernelChannel_CP_676_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_349/do_while_stmt_350/loop_back
      -- 
    -- Element group loadKernelChannel_CP_676_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	88 
    -- CP-element group 14: 	89 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/condition_done
      -- 
    loadKernelChannel_CP_676_elements(14) <= loadKernelChannel_CP_676_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	87 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_349/do_while_stmt_350/loop_body_done
      -- 
    loadKernelChannel_CP_676_elements(15) <= loadKernelChannel_CP_676_elements(87);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_676_elements(16) <= loadKernelChannel_CP_676_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_676_elements(17) <= loadKernelChannel_CP_676_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	64 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	86 
    -- CP-element group 18: 	24 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	27 
    -- CP-element group 19: 	86 
    -- CP-element group 19: 	23 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/condition_evaluated
      -- 
    condition_evaluated_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(19), ack => do_while_stmt_350_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(27) & loadKernelChannel_CP_676_elements(86) & loadKernelChannel_CP_676_elements(23);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	41 
    -- CP-element group 20: 	24 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_req
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start__ps
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(41) & loadKernelChannel_CP_676_elements(24) & loadKernelChannel_CP_676_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	75 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	83 
    -- CP-element group 21: 	87 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	41 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(26) & loadKernelChannel_CP_676_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_req
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start__ps
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(25) & loadKernelChannel_CP_676_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(27) & loadKernelChannel_CP_676_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	66 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	80 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(27) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(72) & loadKernelChannel_CP_676_elements(80);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	60 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	70 
    -- CP-element group 27: 	78 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed__ps
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(27), ack => array_obj_ref_397_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(28) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req_ps
      -- 
    phi_stmt_352_loopback_sample_req_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_loopback_sample_req_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(29), ack => phi_stmt_352_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(30) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req
      -- CP-element group 31: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req_ps
      -- 
    phi_stmt_352_entry_sample_req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_entry_sample_req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(31), ack => phi_stmt_352_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack
      -- CP-element group 32: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack_ps
      -- 
    phi_stmt_352_phi_mux_ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_352_ack_0, ack => loadKernelChannel_CP_676_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/req
      -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(33), ack => nmycount_374_354_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start_
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/req
      -- 
    req_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(34), ack => nmycount_374_354_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/ack
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_0, ack => loadKernelChannel_CP_676_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/ack
      -- 
    ack_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_1, ack => loadKernelChannel_CP_676_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start__ps
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/req
      -- 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(37), ack => start_add_355_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start_
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/req
      -- 
    req_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(38), ack => start_add_355_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/ack
      -- 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_0, ack => loadKernelChannel_CP_676_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/ack
      -- 
    ack_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_1, ack => loadKernelChannel_CP_676_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	81 
    -- CP-element group 41: 	85 
    -- CP-element group 41: 	21 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	84 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start__ps
      -- 
    loadKernelChannel_CP_676_elements(43) <= loadKernelChannel_CP_676_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start__ps
      -- 
    loadKernelChannel_CP_676_elements(45) <= loadKernelChannel_CP_676_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	82 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_676_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(47) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req_ps
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req
      -- 
    phi_stmt_356_loopback_sample_req_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_loopback_sample_req_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(48), ack => phi_stmt_356_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(49) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req_ps
      -- 
    phi_stmt_356_entry_sample_req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_entry_sample_req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(50), ack => phi_stmt_356_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack_ps
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack
      -- 
    phi_stmt_356_phi_mux_ack_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_356_ack_0, ack => loadKernelChannel_CP_676_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/req
      -- 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(52), ack => nfetch_val_419_358_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start_
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/req
      -- 
    req_906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(53), ack => nfetch_val_419_358_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$exit
      -- 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_0, ack => loadKernelChannel_CP_676_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/ack
      -- 
    ack_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_1, ack => loadKernelChannel_CP_676_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start_
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(56), ack => my_fetch_339_359_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start_
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/req
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start__ps
      -- 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(57), ack => my_fetch_339_359_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed__ps
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_0, ack => loadKernelChannel_CP_676_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed__ps
      -- 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_1, ack => loadKernelChannel_CP_676_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/req
      -- 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(60), ack => WPIPE_kernel_pipe1_381_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(27) & loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_start_
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/req
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$exit
      -- 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_0, ack => loadKernelChannel_CP_676_elements(61)); -- 
    req_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(61), ack => WPIPE_kernel_pipe1_381_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	87 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$exit
      -- 
    ack_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_1, ack => loadKernelChannel_CP_676_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	67 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	68 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$entry
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/req
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_start_
      -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(63), ack => addr_of_398_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	18 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: 	76 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/req
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_start_
      -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(64), ack => addr_of_398_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(69) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_update_start
      -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(65), ack => array_obj_ref_397_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	25 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_sample_complete
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (8) 
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_offset_calculated
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_req
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_root_address_calculated
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	65 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$exit
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/ack
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_completed_
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	64 
    -- CP-element group 69:  members (19) 
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_root_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_resized
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_req
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	27 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(70), ack => W_fn_388_delayed_7_0_400_inst_req_0); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(27) & loadKernelChannel_CP_676_elements(72);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	76 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/req
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_start_
      -- 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(71), ack => W_fn_388_delayed_7_0_400_inst_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	25 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/ack
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_0, ack => loadKernelChannel_CP_676_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_completed_
      -- 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_1, ack => loadKernelChannel_CP_676_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	73 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/rr
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$entry
      -- 
    rr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(74), ack => ptr_deref_406_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(69) & loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	21 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_start_
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$entry
      -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(75), ack => ptr_deref_406_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(77);
      gj_loadKernelChannel_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	64 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/ra
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$exit
      -- 
    ra_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	87 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_ack
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_req
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$entry
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/ca
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$exit
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	27 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/req
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_start_
      -- 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(78), ack => W_fn_394_delayed_13_0_408_inst_req_0); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(27) & loadKernelChannel_CP_676_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	21 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_start_
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/req
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$entry
      -- 
    req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(79), ack => W_fn_394_delayed_13_0_408_inst_req_1); -- 
    loadKernelChannel_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(81);
      gj_loadKernelChannel_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	25 
    -- CP-element group 80: 	78 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/ack
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_completed_
      -- 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_0, ack => loadKernelChannel_CP_676_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	41 
    -- CP-element group 81: 	79 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/ack
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$exit
      -- 
    ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_1, ack => loadKernelChannel_CP_676_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	46 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/req
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(82), ack => W_fetch_val_396_delayed_13_0_411_inst_req_0); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	21 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/req
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_start_
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$entry
      -- 
    req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(83), ack => W_fetch_val_396_delayed_13_0_411_inst_req_1); -- 
    loadKernelChannel_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(85);
      gj_loadKernelChannel_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	42 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/ack
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_completed_
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_0, ack => loadKernelChannel_CP_676_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	41 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_completed_
      -- 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_1, ack => loadKernelChannel_CP_676_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	18 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	19 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_676_elements(18), ack => loadKernelChannel_CP_676_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	62 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	77 
    -- CP-element group 87: 	81 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	21 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	15 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(62) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	14 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$exit
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/ack
      -- 
    ack_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_0, ack => loadKernelChannel_CP_676_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	14 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/ack
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$exit
      -- 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_1, ack => loadKernelChannel_CP_676_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	12 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	10 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_349/do_while_stmt_350/$exit
      -- 
    loadKernelChannel_CP_676_elements(90) <= loadKernelChannel_CP_676_elements(12);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	10 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_sample_completed_
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/$exit
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/ra
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_0, ack => loadKernelChannel_CP_676_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	10 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/req
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_start_
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/ca
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_update_completed_
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/$exit
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_1, ack => loadKernelChannel_CP_676_elements(92)); -- 
    req_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(92), ack => WPIPE_size_pipe_428_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_completed_
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/ack
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/req
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$exit
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$entry
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_update_start_
      -- 
    ack_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_0, ack => loadKernelChannel_CP_676_elements(93)); -- 
    req_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(93), ack => WPIPE_size_pipe_428_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 assign_stmt_433/$exit
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_update_completed_
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$exit
      -- CP-element group 94: 	 $exit
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/ack
      -- 
    ack_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_1, ack => loadKernelChannel_CP_676_elements(94)); -- 
    loadKernelChannel_do_while_stmt_350_terminator_1088: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_350_terminator_1088", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_676_elements(15),loop_continue => loadKernelChannel_CP_676_elements(89),loop_terminate => loadKernelChannel_CP_676_elements(88),loop_back => loadKernelChannel_CP_676_elements(13),loop_exit => loadKernelChannel_CP_676_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_352_phi_seq_872_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(28);
      loadKernelChannel_CP_676_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(35);
      loadKernelChannel_CP_676_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(36);
      loadKernelChannel_CP_676_elements(29) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(30);
      loadKernelChannel_CP_676_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(39);
      loadKernelChannel_CP_676_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(40);
      loadKernelChannel_CP_676_elements(31) <= phi_mux_reqs(1);
      phi_stmt_352_phi_seq_872 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_352_phi_seq_872") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(26), 
          phi_update_req => loadKernelChannel_CP_676_elements(22), 
          phi_update_ack => loadKernelChannel_CP_676_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_356_phi_seq_926_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(47);
      loadKernelChannel_CP_676_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(54);
      loadKernelChannel_CP_676_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(55);
      loadKernelChannel_CP_676_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(49);
      loadKernelChannel_CP_676_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(58);
      loadKernelChannel_CP_676_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(59);
      loadKernelChannel_CP_676_elements(50) <= phi_mux_reqs(1);
      phi_stmt_356_phi_seq_926 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_356_phi_seq_926") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(44), 
          phi_update_req => loadKernelChannel_CP_676_elements(45), 
          phi_update_ack => loadKernelChannel_CP_676_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_814_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_676_elements(16);
        preds(1)  <= loadKernelChannel_CP_676_elements(17);
        entry_tmerge_814 : transition_merge -- 
          generic map(name => " entry_tmerge_814")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_676_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_365_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_387_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_378_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_396_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_332_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_332_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_366_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_424_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_431_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_425_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_333_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_335 : std_logic_vector(31 downto 0);
    signal fetch_addr_399 : std_logic_vector(31 downto 0);
    signal fetch_val_356 : std_logic_vector(63 downto 0);
    signal fetch_val_396_delayed_13_0_413 : std_logic_vector(63 downto 0);
    signal first_fill_344 : std_logic_vector(0 downto 0);
    signal fn_388_delayed_7_0_402 : std_logic_vector(0 downto 0);
    signal fn_390 : std_logic_vector(0 downto 0);
    signal fn_394_delayed_13_0_410 : std_logic_vector(0 downto 0);
    signal fv_407 : std_logic_vector(63 downto 0);
    signal konst_326_wire_constant : std_logic_vector(63 downto 0);
    signal konst_342_wire_constant : std_logic_vector(63 downto 0);
    signal konst_362_wire_constant : std_logic_vector(63 downto 0);
    signal konst_364_wire_constant : std_logic_vector(63 downto 0);
    signal konst_367_wire_constant : std_logic_vector(63 downto 0);
    signal konst_372_wire_constant : std_logic_vector(63 downto 0);
    signal konst_386_wire_constant : std_logic_vector(63 downto 0);
    signal konst_388_wire_constant : std_logic_vector(63 downto 0);
    signal konst_395_wire_constant : std_logic_vector(63 downto 0);
    signal konst_423_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_339 : std_logic_vector(63 downto 0);
    signal my_fetch_339_359_buffered : std_logic_vector(63 downto 0);
    signal my_num1_369 : std_logic_vector(63 downto 0);
    signal mycount_352 : std_logic_vector(63 downto 0);
    signal nfetch_val_419 : std_logic_vector(63 downto 0);
    signal nfetch_val_419_358_buffered : std_logic_vector(63 downto 0);
    signal nmycount_374 : std_logic_vector(63 downto 0);
    signal nmycount_374_354_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_338_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_338_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_406_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_328 : std_logic_vector(63 downto 0);
    signal start_add_355_buffered : std_logic_vector(63 downto 0);
    signal start_next_348 : std_logic_vector(0 downto 0);
    signal type_cast_432_wire : std_logic_vector(31 downto 0);
    signal var_val_380 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_333_constant_part_of_offset <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_333_resized_base_address <= "00000000000000";
    array_obj_ref_397_constant_part_of_offset <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_397_resized_base_address <= "00000000000000";
    konst_326_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_362_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_367_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_372_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_388_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_395_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_338_word_offset_0 <= "00000000000000";
    ptr_deref_406_word_offset_0 <= "00000000000000";
    phi_stmt_352: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_374_354_buffered & start_add_355_buffered;
      req <= phi_stmt_352_req_0 & phi_stmt_352_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_352",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_352_ack_0,
          idata => idata,
          odata => mycount_352,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_352
    phi_stmt_356: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_419_358_buffered & my_fetch_339_359_buffered;
      req <= phi_stmt_356_req_0 & phi_stmt_356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_356",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_356_ack_0,
          idata => idata,
          odata => fetch_val_356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_356
    -- flow-through select operator MUX_418_inst
    nfetch_val_419 <= fv_407 when (fn_394_delayed_13_0_410(0) /=  '0') else fetch_val_396_delayed_13_0_413;
    W_fetch_val_396_delayed_13_0_411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_0;
      W_fetch_val_396_delayed_13_0_411_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_1;
      W_fetch_val_396_delayed_13_0_411_inst_ack_1<= rack(0);
      W_fetch_val_396_delayed_13_0_411_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_396_delayed_13_0_411_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_396_delayed_13_0_413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_388_delayed_7_0_400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_388_delayed_7_0_400_inst_req_0;
      W_fn_388_delayed_7_0_400_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_388_delayed_7_0_400_inst_req_1;
      W_fn_388_delayed_7_0_400_inst_ack_1<= rack(0);
      W_fn_388_delayed_7_0_400_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_388_delayed_7_0_400_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_388_delayed_7_0_402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_394_delayed_13_0_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_394_delayed_13_0_408_inst_req_0;
      W_fn_394_delayed_13_0_408_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_394_delayed_13_0_408_inst_req_1;
      W_fn_394_delayed_13_0_408_inst_ack_1<= rack(0);
      W_fn_394_delayed_13_0_408_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_394_delayed_13_0_408_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_394_delayed_13_0_410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_334_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_334_final_reg_req_0;
      addr_of_334_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_334_final_reg_req_1;
      addr_of_334_final_reg_ack_1<= rack(0);
      addr_of_334_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_334_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_333_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_398_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_398_final_reg_req_0;
      addr_of_398_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_398_final_reg_req_1;
      addr_of_398_final_reg_ack_1<= rack(0);
      addr_of_398_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_398_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_397_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_339_359_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_339_359_buf_req_0;
      my_fetch_339_359_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_339_359_buf_req_1;
      my_fetch_339_359_buf_ack_1<= rack(0);
      my_fetch_339_359_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_339_359_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_339_359_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_419_358_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_419_358_buf_req_0;
      nfetch_val_419_358_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_419_358_buf_req_1;
      nfetch_val_419_358_buf_ack_1<= rack(0);
      nfetch_val_419_358_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_419_358_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_419_358_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_374_354_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_374_354_buf_req_0;
      nmycount_374_354_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_374_354_buf_req_1;
      nmycount_374_354_buf_ack_1<= rack(0);
      nmycount_374_354_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_374_354_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_374_354_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_355_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_355_buf_req_0;
      start_add_355_buf_ack_0<= wack(0);
      rreq(0) <= start_add_355_buf_req_1;
      start_add_355_buf_ack_1<= rack(0);
      start_add_355_buf : InterlockBuffer generic map ( -- 
        name => "start_add_355_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_355_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_379_inst
    process(LSHR_u64_u64_378_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_378_wire(15 downto 0);
      var_val_380 <= tmp_var; -- 
    end process;
    type_cast_432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_432_inst_req_0;
      type_cast_432_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_432_inst_req_1;
      type_cast_432_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  first_fill_344(0);
      type_cast_432_inst_gI: SplitGuardInterface generic map(name => "type_cast_432_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SUB_u64_u64_431_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_333_index_1_rename
    process(R_sh_start_332_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_332_resized;
      ov(13 downto 0) := iv;
      R_sh_start_332_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_index_1_resize
    process(sh_start_328) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_328;
      ov := iv(13 downto 0);
      R_sh_start_332_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_root_address_inst
    process(array_obj_ref_333_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_333_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_333_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_rename
    process(LSHR_u64_u64_396_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_396_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_resize
    process(LSHR_u64_u64_396_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_396_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_root_address_inst
    process(array_obj_ref_397_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_397_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_397_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_addr_0
    process(ptr_deref_338_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_base_resize
    process(fetch_addr_335) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_335;
      ov := iv(13 downto 0);
      ptr_deref_338_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_gather_scatter
    process(ptr_deref_338_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_data_0;
      ov(63 downto 0) := iv;
      my_fetch_339 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_root_address_inst
    process(ptr_deref_338_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_addr_0
    process(ptr_deref_406_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_base_resize
    process(fetch_addr_399) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_399;
      ov := iv(13 downto 0);
      ptr_deref_406_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_gather_scatter
    process(ptr_deref_406_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_data_0;
      ov(63 downto 0) := iv;
      fv_407 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_root_address_inst
    process(ptr_deref_406_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_350_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_425_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_350_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_350_branch_req_0,
          ack0 => do_while_stmt_350_branch_ack_0,
          ack1 => do_while_stmt_350_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_373_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_352, konst_372_wire_constant, tmp_var);
      nmycount_374 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_365_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_352, konst_364_wire_constant, tmp_var);
      AND_u64_u64_365_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_387_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_374, konst_386_wire_constant, tmp_var);
      AND_u64_u64_387_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_343_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_342_wire_constant, tmp_var);
      first_fill_344 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_389_inst
    process(AND_u64_u64_387_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_387_wire, konst_388_wire_constant, tmp_var);
      fn_390 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_327_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_326_wire_constant, tmp_var);
      sh_start_328 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_378_inst
    process(fetch_val_356, my_num1_369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_356, my_num1_369, tmp_var);
      LSHR_u64_u64_378_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_396_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_374, konst_395_wire_constant, tmp_var);
      LSHR_u64_u64_396_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_368_inst
    process(SUB_u64_u64_366_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_366_wire, konst_367_wire_constant, tmp_var);
      my_num1_369 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_366_inst
    process(konst_362_wire_constant, AND_u64_u64_365_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_362_wire_constant, AND_u64_u64_365_wire, tmp_var);
      SUB_u64_u64_366_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_424_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_423_wire_constant, tmp_var);
      SUB_u64_u64_424_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_431_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_431_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_425_inst
    process(mycount_352, SUB_u64_u64_424_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_352, SUB_u64_u64_424_wire, tmp_var);
      ULT_u64_u1_425_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : array_obj_ref_333_index_offset 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_332_scaled;
      array_obj_ref_333_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_333_index_offset_req_0;
      array_obj_ref_333_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_333_index_offset_req_1;
      array_obj_ref_333_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_397_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_396_scaled;
      array_obj_ref_397_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_397_index_offset_req_0;
      array_obj_ref_397_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_397_index_offset_req_1;
      array_obj_ref_397_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_338_load_0 ptr_deref_406_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_338_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_406_load_0_req_0;
      ptr_deref_338_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_406_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_338_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_406_load_0_req_1;
      ptr_deref_338_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_406_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_388_delayed_7_0_402(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_338_word_address_0 & ptr_deref_406_word_address_0;
      ptr_deref_338_data_0 <= data_out(127 downto 64);
      ptr_deref_406_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_347_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_0;
      RPIPE_input_done_pipe_347_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_1;
      RPIPE_input_done_pipe_347_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_344(0);
      start_next_348 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_381_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_0;
      WPIPE_kernel_pipe1_381_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_1;
      WPIPE_kernel_pipe1_381_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val_380;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_size_pipe_428_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_0;
      WPIPE_size_pipe_428_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_1;
      WPIPE_size_pipe_428_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= first_fill_344(0);
      data_in <= type_cast_432_wire;
      size_pipe_write_1_gI: SplitGuardInterface generic map(name => "size_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_318_load_0_req_0 : boolean;
  signal LOAD_count_318_load_0_ack_0 : boolean;
  signal LOAD_count_318_load_0_req_1 : boolean;
  signal LOAD_count_318_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_319/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_sample_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_update_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/cr
      -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_1); -- 
    rr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_sample_completed_
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/ra
      -- 
    ra_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_0, ack => timer_CP_637_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_319/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_update_completed_
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_ack
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_1, ack => timer_CP_637_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_318_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_318_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_318_word_address_0 <= "0";
    -- equivalence LOAD_count_318_gather_scatter
    process(LOAD_count_318_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_318_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_318_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_318_load_0_req_0;
      LOAD_count_318_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_318_load_0_req_1;
      LOAD_count_318_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_318_word_address_0;
      LOAD_count_318_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_4562_start: Boolean;
  signal timerDaemon_CP_4562_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1997_branch_req_0 : boolean;
  signal phi_stmt_1999_req_0 : boolean;
  signal phi_stmt_1999_req_1 : boolean;
  signal phi_stmt_1999_ack_0 : boolean;
  signal ADD_u64_u64_2003_inst_req_0 : boolean;
  signal ADD_u64_u64_2003_inst_ack_0 : boolean;
  signal ADD_u64_u64_2003_inst_req_1 : boolean;
  signal ADD_u64_u64_2003_inst_ack_1 : boolean;
  signal STORE_count_2007_store_0_req_0 : boolean;
  signal STORE_count_2007_store_0_ack_0 : boolean;
  signal STORE_count_2007_store_0_req_1 : boolean;
  signal STORE_count_2007_store_0_ack_1 : boolean;
  signal do_while_stmt_1997_branch_ack_0 : boolean;
  signal do_while_stmt_1997_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_4562_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4562_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_4562_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4562_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_4562: Block -- control-path 
    signal timerDaemon_CP_4562_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_4562_elements(0) <= timerDaemon_CP_4562_start;
    timerDaemon_CP_4562_symbol <= timerDaemon_CP_4562_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1996/$entry
      -- CP-element group 0: 	 branch_block_stmt_1996/branch_block_stmt_1996__entry__
      -- CP-element group 0: 	 branch_block_stmt_1996/do_while_stmt_1997__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1996/$exit
      -- CP-element group 1: 	 branch_block_stmt_1996/branch_block_stmt_1996__exit__
      -- CP-element group 1: 	 branch_block_stmt_1996/do_while_stmt_1997__exit__
      -- 
    timerDaemon_CP_4562_elements(1) <= timerDaemon_CP_4562_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1996/do_while_stmt_1997/$entry
      -- CP-element group 2: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997__entry__
      -- 
    timerDaemon_CP_4562_elements(2) <= timerDaemon_CP_4562_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997__exit__
      -- 
    -- Element group timerDaemon_CP_4562_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_back
      -- 
    -- Element group timerDaemon_CP_4562_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1996/do_while_stmt_1997/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_taken/$entry
      -- 
    timerDaemon_CP_4562_elements(5) <= timerDaemon_CP_4562_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_body_done
      -- 
    timerDaemon_CP_4562_elements(6) <= timerDaemon_CP_4562_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_4562_elements(7) <= timerDaemon_CP_4562_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_4562_elements(8) <= timerDaemon_CP_4562_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_4562_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/condition_evaluated
      -- 
    condition_evaluated_4586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4562_elements(10), ack => do_while_stmt_1997_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(35) & timerDaemon_CP_4562_elements(15);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(12) & timerDaemon_CP_4562_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(9) & timerDaemon_CP_4562_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(9) & timerDaemon_CP_4562_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_4562_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_4562_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_loopback_trigger
      -- 
    timerDaemon_CP_4562_elements(16) <= timerDaemon_CP_4562_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_loopback_sample_req_ps
      -- 
    phi_stmt_1999_loopback_sample_req_4601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1999_loopback_sample_req_4601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4562_elements(17), ack => phi_stmt_1999_req_0); -- 
    -- Element group timerDaemon_CP_4562_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_entry_trigger
      -- 
    timerDaemon_CP_4562_elements(18) <= timerDaemon_CP_4562_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_entry_sample_req_ps
      -- 
    phi_stmt_1999_entry_sample_req_4604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1999_entry_sample_req_4604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4562_elements(19), ack => phi_stmt_1999_req_1); -- 
    -- Element group timerDaemon_CP_4562_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/phi_stmt_1999_phi_mux_ack_ps
      -- 
    phi_stmt_1999_phi_mux_ack_4607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1999_ack_0, ack => timerDaemon_CP_4562_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_4562_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_update_start__ps
      -- 
    -- Element group timerDaemon_CP_4562_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Sample/rr
      -- 
    rr_4620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4562_elements(23), ack => ADD_u64_u64_2003_inst_req_0); -- 
    timerDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(21) & timerDaemon_CP_4562_elements(25);
      gj_timerDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Update/cr
      -- 
    cr_4625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4562_elements(24), ack => ADD_u64_u64_2003_inst_req_1); -- 
    timerDaemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(22) & timerDaemon_CP_4562_elements(26);
      gj_timerDaemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Sample/ra
      -- 
    ra_4621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2003_inst_ack_0, ack => timerDaemon_CP_4562_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_update_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/ADD_u64_u64_2003_Update/ca
      -- 
    ca_4626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2003_inst_ack_1, ack => timerDaemon_CP_4562_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_sample_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_sample_completed_
      -- 
    -- Element group timerDaemon_CP_4562_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_update_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_update_start_
      -- 
    -- Element group timerDaemon_CP_4562_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_update_completed__ps
      -- 
    timerDaemon_CP_4562_elements(29) <= timerDaemon_CP_4562_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/type_cast_2005_update_completed_
      -- 
    -- Element group timerDaemon_CP_4562_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => timerDaemon_CP_4562_elements(28), ack => timerDaemon_CP_4562_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/STORE_count_2007_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/STORE_count_2007_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/STORE_count_2007_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/STORE_count_2007_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/word_access_start/word_0/rr
      -- 
    rr_4656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4562_elements(31), ack => STORE_count_2007_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(9) & timerDaemon_CP_4562_elements(15) & timerDaemon_CP_4562_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/word_access_complete/word_0/cr
      -- 
    cr_4667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4562_elements(32), ack => STORE_count_2007_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_4562_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Sample/word_access_start/word_0/ra
      -- 
    ra_4657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2007_store_0_ack_0, ack => timerDaemon_CP_4562_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/STORE_count_2007_Update/word_access_complete/word_0/ca
      -- 
    ca_4668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2007_store_0_ack_1, ack => timerDaemon_CP_4562_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_4562_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_4562_elements(9), ack => timerDaemon_CP_4562_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1996/do_while_stmt_1997/do_while_stmt_1997_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4562_elements(14) & timerDaemon_CP_4562_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4562_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_exit/ack
      -- 
    ack_4673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1997_branch_ack_0, ack => timerDaemon_CP_4562_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_1996/do_while_stmt_1997/loop_taken/ack
      -- 
    ack_4677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1997_branch_ack_1, ack => timerDaemon_CP_4562_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1996/do_while_stmt_1997/$exit
      -- 
    timerDaemon_CP_4562_elements(39) <= timerDaemon_CP_4562_elements(3);
    timerDaemon_do_while_stmt_1997_terminator_4678: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1997_terminator_4678", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_4562_elements(6),loop_continue => timerDaemon_CP_4562_elements(38),loop_terminate => timerDaemon_CP_4562_elements(37),loop_back => timerDaemon_CP_4562_elements(4),loop_exit => timerDaemon_CP_4562_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1999_phi_seq_4635_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_4562_elements(16);
      timerDaemon_CP_4562_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_4562_elements(25);
      timerDaemon_CP_4562_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_4562_elements(26);
      timerDaemon_CP_4562_elements(17) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_4562_elements(18);
      timerDaemon_CP_4562_elements(27)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_4562_elements(27);
      timerDaemon_CP_4562_elements(28)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_4562_elements(29);
      timerDaemon_CP_4562_elements(19) <= phi_mux_reqs(1);
      phi_stmt_1999_phi_seq_4635 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_1999_phi_seq_4635") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_4562_elements(11), 
          phi_sample_ack => timerDaemon_CP_4562_elements(14), 
          phi_update_req => timerDaemon_CP_4562_elements(13), 
          phi_update_ack => timerDaemon_CP_4562_elements(15), 
          phi_mux_ack => timerDaemon_CP_4562_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4587_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_4562_elements(7);
        preds(1)  <= timerDaemon_CP_4562_elements(8);
        entry_tmerge_4587 : transition_merge -- 
          generic map(name => " entry_tmerge_4587")
          port map (preds => preds, symbol_out => timerDaemon_CP_4562_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_2003_wire : std_logic_vector(63 downto 0);
    signal STORE_count_2007_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_2007_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_2002_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2011_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_1999 : std_logic_vector(63 downto 0);
    signal type_cast_2005_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_2007_word_address_0 <= "0";
    konst_2002_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2011_wire_constant <= "1";
    type_cast_2005_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1999: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u64_u64_2003_wire & type_cast_2005_wire_constant;
      req <= phi_stmt_1999_req_0 & phi_stmt_1999_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1999",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1999_ack_0,
          idata => idata,
          odata => ncount_1999,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1999
    -- equivalence STORE_count_2007_gather_scatter
    process(ncount_1999) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_1999;
      ov(63 downto 0) := iv;
      STORE_count_2007_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_1997_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2011_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1997_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1997_branch_req_0,
          ack0 => do_while_stmt_1997_branch_ack_0,
          ack1 => do_while_stmt_1997_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_2003_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_1999;
      ADD_u64_u64_2003_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2003_inst_req_0;
      ADD_u64_u64_2003_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2003_inst_req_1;
      ADD_u64_u64_2003_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_2007_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_2007_store_0_req_0;
      STORE_count_2007_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_2007_store_0_req_1;
      STORE_count_2007_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_2007_word_address_0;
      data_in <= STORE_count_2007_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(127 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(127 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(127 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(127 downto 64);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(63 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 128,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
