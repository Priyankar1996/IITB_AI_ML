-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    row_in : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal row_in_buffer :  std_logic_vector(15 downto 0);
  signal row_in_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_359_load_0_ack_1 : boolean;
  signal ptr_deref_359_load_0_req_1 : boolean;
  signal W_fn2_265_delayed_13_0_282_inst_req_0 : boolean;
  signal addr_of_272_final_reg_ack_0 : boolean;
  signal addr_of_272_final_reg_req_0 : boolean;
  signal W_fn2_259_delayed_7_0_274_inst_ack_1 : boolean;
  signal W_fn2_259_delayed_7_0_274_inst_req_1 : boolean;
  signal ptr_deref_51_load_0_req_0 : boolean;
  signal ptr_deref_51_load_0_ack_0 : boolean;
  signal ptr_deref_51_load_0_req_1 : boolean;
  signal ptr_deref_51_load_0_ack_1 : boolean;
  signal array_obj_ref_74_index_offset_req_0 : boolean;
  signal array_obj_ref_74_index_offset_ack_0 : boolean;
  signal array_obj_ref_60_index_offset_req_0 : boolean;
  signal array_obj_ref_60_index_offset_ack_0 : boolean;
  signal array_obj_ref_60_index_offset_req_1 : boolean;
  signal array_obj_ref_60_index_offset_ack_1 : boolean;
  signal WPIPE_input_pipe2_294_inst_ack_1 : boolean;
  signal ptr_deref_280_load_0_ack_0 : boolean;
  signal array_obj_ref_350_index_offset_ack_0 : boolean;
  signal addr_of_61_final_reg_req_0 : boolean;
  signal addr_of_61_final_reg_ack_0 : boolean;
  signal addr_of_61_final_reg_req_1 : boolean;
  signal addr_of_61_final_reg_ack_1 : boolean;
  signal ptr_deref_280_load_0_req_0 : boolean;
  signal W_fn2_259_delayed_7_0_274_inst_ack_0 : boolean;
  signal W_fn2_259_delayed_7_0_274_inst_req_0 : boolean;
  signal ptr_deref_65_load_0_req_0 : boolean;
  signal ptr_deref_65_load_0_ack_0 : boolean;
  signal ptr_deref_65_load_0_req_1 : boolean;
  signal ptr_deref_65_load_0_ack_1 : boolean;
  signal WPIPE_input_pipe2_294_inst_req_1 : boolean;
  signal ptr_deref_280_load_0_ack_1 : boolean;
  signal addr_of_351_final_reg_ack_1 : boolean;
  signal W_fn3_332_delayed_13_0_361_inst_req_1 : boolean;
  signal W_fn3_332_delayed_13_0_361_inst_ack_1 : boolean;
  signal W_fn3_326_delayed_7_0_353_inst_ack_0 : boolean;
  signal W_fn3_326_delayed_7_0_353_inst_req_0 : boolean;
  signal array_obj_ref_350_index_offset_req_0 : boolean;
  signal array_obj_ref_74_index_offset_req_1 : boolean;
  signal array_obj_ref_74_index_offset_ack_1 : boolean;
  signal addr_of_75_final_reg_req_0 : boolean;
  signal addr_of_75_final_reg_ack_0 : boolean;
  signal addr_of_75_final_reg_req_1 : boolean;
  signal addr_of_75_final_reg_ack_1 : boolean;
  signal W_continue_247_delayed_1_0_251_inst_ack_1 : boolean;
  signal ptr_deref_280_load_0_req_1 : boolean;
  signal ptr_deref_79_load_0_req_0 : boolean;
  signal ptr_deref_79_load_0_ack_0 : boolean;
  signal ptr_deref_79_load_0_req_1 : boolean;
  signal ptr_deref_79_load_0_ack_1 : boolean;
  signal addr_of_351_final_reg_req_1 : boolean;
  signal array_obj_ref_271_index_offset_ack_1 : boolean;
  signal do_while_stmt_81_branch_req_0 : boolean;
  signal array_obj_ref_271_index_offset_req_1 : boolean;
  signal W_fetch_val2_267_delayed_13_0_285_inst_ack_1 : boolean;
  signal WPIPE_input_pipe2_294_inst_ack_0 : boolean;
  signal W_fetch_val2_267_delayed_13_0_285_inst_req_1 : boolean;
  signal phi_stmt_83_req_1 : boolean;
  signal W_fn3_332_delayed_13_0_361_inst_req_0 : boolean;
  signal phi_stmt_83_req_0 : boolean;
  signal phi_stmt_83_ack_0 : boolean;
  signal WPIPE_input_pipe2_294_inst_req_0 : boolean;
  signal W_fetch_val2_267_delayed_13_0_285_inst_ack_0 : boolean;
  signal W_fn3_326_delayed_7_0_353_inst_ack_1 : boolean;
  signal W_fetch_val2_267_delayed_13_0_285_inst_req_0 : boolean;
  signal n_address1_176_87_buf_req_0 : boolean;
  signal n_address1_176_87_buf_ack_0 : boolean;
  signal array_obj_ref_271_index_offset_ack_0 : boolean;
  signal W_continue_309_delayed_1_0_325_inst_ack_1 : boolean;
  signal n_address1_176_87_buf_req_1 : boolean;
  signal n_address1_176_87_buf_ack_1 : boolean;
  signal W_fn3_326_delayed_7_0_353_inst_req_1 : boolean;
  signal addr_of_272_final_reg_ack_1 : boolean;
  signal W_continue_309_delayed_1_0_325_inst_req_1 : boolean;
  signal phi_stmt_88_req_1 : boolean;
  signal phi_stmt_88_req_0 : boolean;
  signal W_continue_309_delayed_1_0_325_inst_ack_0 : boolean;
  signal array_obj_ref_271_index_offset_req_0 : boolean;
  signal phi_stmt_88_ack_0 : boolean;
  signal addr_of_351_final_reg_ack_0 : boolean;
  signal W_continue_309_delayed_1_0_325_inst_req_0 : boolean;
  signal type_cast_91_inst_req_0 : boolean;
  signal type_cast_91_inst_ack_0 : boolean;
  signal type_cast_91_inst_req_1 : boolean;
  signal type_cast_91_inst_ack_1 : boolean;
  signal phi_stmt_115_req_1 : boolean;
  signal phi_stmt_115_req_0 : boolean;
  signal phi_stmt_115_ack_0 : boolean;
  signal n_address2_250_92_buf_req_0 : boolean;
  signal n_address2_250_92_buf_ack_0 : boolean;
  signal n_address2_250_92_buf_req_1 : boolean;
  signal n_address2_250_92_buf_ack_1 : boolean;
  signal addr_of_272_final_reg_req_1 : boolean;
  signal ptr_deref_359_load_0_ack_0 : boolean;
  signal phi_stmt_93_req_1 : boolean;
  signal phi_stmt_93_req_0 : boolean;
  signal phi_stmt_93_ack_0 : boolean;
  signal addr_of_351_final_reg_req_0 : boolean;
  signal type_cast_96_inst_req_0 : boolean;
  signal type_cast_96_inst_ack_0 : boolean;
  signal type_cast_96_inst_req_1 : boolean;
  signal type_cast_96_inst_ack_1 : boolean;
  signal array_obj_ref_350_index_offset_ack_1 : boolean;
  signal ptr_deref_359_load_0_req_0 : boolean;
  signal n_address3_324_97_buf_req_0 : boolean;
  signal n_address3_324_97_buf_ack_0 : boolean;
  signal n_address3_324_97_buf_req_1 : boolean;
  signal n_address3_324_97_buf_ack_1 : boolean;
  signal array_obj_ref_350_index_offset_req_1 : boolean;
  signal phi_stmt_98_req_1 : boolean;
  signal W_fn3_332_delayed_13_0_361_inst_ack_0 : boolean;
  signal phi_stmt_98_req_0 : boolean;
  signal phi_stmt_98_ack_0 : boolean;
  signal W_fn2_265_delayed_13_0_282_inst_ack_1 : boolean;
  signal W_fn2_265_delayed_13_0_282_inst_req_1 : boolean;
  signal W_fn2_265_delayed_13_0_282_inst_ack_0 : boolean;
  signal n_mycounter_143_102_buf_req_0 : boolean;
  signal n_mycounter_143_102_buf_ack_0 : boolean;
  signal n_mycounter_143_102_buf_req_1 : boolean;
  signal n_mycounter_143_102_buf_ack_1 : boolean;
  signal phi_stmt_103_req_1 : boolean;
  signal phi_stmt_103_req_0 : boolean;
  signal phi_stmt_103_ack_0 : boolean;
  signal my_fetch1_52_105_buf_req_0 : boolean;
  signal my_fetch1_52_105_buf_ack_0 : boolean;
  signal my_fetch1_52_105_buf_req_1 : boolean;
  signal my_fetch1_52_105_buf_ack_1 : boolean;
  signal W_continue_247_delayed_1_0_251_inst_req_1 : boolean;
  signal n_fetch_val1_219_106_buf_req_0 : boolean;
  signal n_fetch_val1_219_106_buf_ack_0 : boolean;
  signal n_fetch_val1_219_106_buf_req_1 : boolean;
  signal n_fetch_val1_219_106_buf_ack_1 : boolean;
  signal phi_stmt_107_req_1 : boolean;
  signal phi_stmt_107_req_0 : boolean;
  signal phi_stmt_107_ack_0 : boolean;
  signal my_fetch2_66_109_buf_req_0 : boolean;
  signal my_fetch2_66_109_buf_ack_0 : boolean;
  signal my_fetch2_66_109_buf_req_1 : boolean;
  signal my_fetch2_66_109_buf_ack_1 : boolean;
  signal n_fetch_val2_293_110_buf_req_0 : boolean;
  signal n_fetch_val2_293_110_buf_ack_0 : boolean;
  signal n_fetch_val2_293_110_buf_req_1 : boolean;
  signal n_fetch_val2_293_110_buf_ack_1 : boolean;
  signal phi_stmt_111_req_1 : boolean;
  signal phi_stmt_111_req_0 : boolean;
  signal phi_stmt_111_ack_0 : boolean;
  signal my_fetch3_80_113_buf_req_0 : boolean;
  signal my_fetch3_80_113_buf_ack_0 : boolean;
  signal my_fetch3_80_113_buf_req_1 : boolean;
  signal my_fetch3_80_113_buf_ack_1 : boolean;
  signal n_fetch_val3_372_114_buf_req_0 : boolean;
  signal n_fetch_val3_372_114_buf_ack_0 : boolean;
  signal n_fetch_val3_372_114_buf_req_1 : boolean;
  signal n_fetch_val3_372_114_buf_ack_1 : boolean;
  signal n_row1_171_119_buf_req_0 : boolean;
  signal n_row1_171_119_buf_ack_0 : boolean;
  signal n_row1_171_119_buf_req_1 : boolean;
  signal n_row1_171_119_buf_ack_1 : boolean;
  signal phi_stmt_120_req_1 : boolean;
  signal phi_stmt_120_req_0 : boolean;
  signal phi_stmt_120_ack_0 : boolean;
  signal n_row2_245_124_buf_req_0 : boolean;
  signal n_row2_245_124_buf_ack_0 : boolean;
  signal n_row2_245_124_buf_req_1 : boolean;
  signal n_row2_245_124_buf_ack_1 : boolean;
  signal phi_stmt_125_req_1 : boolean;
  signal phi_stmt_125_req_0 : boolean;
  signal phi_stmt_125_ack_0 : boolean;
  signal n_row3_319_129_buf_req_0 : boolean;
  signal n_row3_319_129_buf_ack_0 : boolean;
  signal n_row3_319_129_buf_req_1 : boolean;
  signal n_row3_319_129_buf_ack_1 : boolean;
  signal W_continue_185_delayed_1_0_177_inst_req_0 : boolean;
  signal W_continue_185_delayed_1_0_177_inst_ack_0 : boolean;
  signal W_continue_185_delayed_1_0_177_inst_req_1 : boolean;
  signal W_continue_185_delayed_1_0_177_inst_ack_1 : boolean;
  signal array_obj_ref_197_index_offset_req_0 : boolean;
  signal array_obj_ref_197_index_offset_ack_0 : boolean;
  signal array_obj_ref_197_index_offset_req_1 : boolean;
  signal array_obj_ref_197_index_offset_ack_1 : boolean;
  signal addr_of_198_final_reg_req_0 : boolean;
  signal addr_of_198_final_reg_ack_0 : boolean;
  signal addr_of_198_final_reg_req_1 : boolean;
  signal addr_of_198_final_reg_ack_1 : boolean;
  signal W_fn1_197_delayed_7_0_200_inst_req_0 : boolean;
  signal W_fn1_197_delayed_7_0_200_inst_ack_0 : boolean;
  signal W_fn1_197_delayed_7_0_200_inst_req_1 : boolean;
  signal W_fn1_197_delayed_7_0_200_inst_ack_1 : boolean;
  signal ptr_deref_206_load_0_req_0 : boolean;
  signal ptr_deref_206_load_0_ack_0 : boolean;
  signal ptr_deref_206_load_0_req_1 : boolean;
  signal ptr_deref_206_load_0_ack_1 : boolean;
  signal W_fn1_203_delayed_13_0_208_inst_req_0 : boolean;
  signal W_fn1_203_delayed_13_0_208_inst_ack_0 : boolean;
  signal W_fn1_203_delayed_13_0_208_inst_req_1 : boolean;
  signal W_fn1_203_delayed_13_0_208_inst_ack_1 : boolean;
  signal W_fetch_val1_205_delayed_13_0_211_inst_req_0 : boolean;
  signal W_fetch_val1_205_delayed_13_0_211_inst_ack_0 : boolean;
  signal W_fetch_val1_205_delayed_13_0_211_inst_req_1 : boolean;
  signal W_fetch_val1_205_delayed_13_0_211_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_220_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_220_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_220_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_220_inst_ack_1 : boolean;
  signal W_continue_247_delayed_1_0_251_inst_req_0 : boolean;
  signal W_continue_247_delayed_1_0_251_inst_ack_0 : boolean;
  signal W_fetch_val3_334_delayed_13_0_364_inst_req_0 : boolean;
  signal W_fetch_val3_334_delayed_13_0_364_inst_ack_0 : boolean;
  signal W_fetch_val3_334_delayed_13_0_364_inst_req_1 : boolean;
  signal W_fetch_val3_334_delayed_13_0_364_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_374_inst_req_0 : boolean;
  signal WPIPE_input_pipe3_374_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_374_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_374_inst_ack_1 : boolean;
  signal do_while_stmt_81_branch_ack_0 : boolean;
  signal do_while_stmt_81_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= row_in;
  row_in_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= ct;
  ct_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(316 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0:  members (79) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_update_start_
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_update_start_
      -- CP-element group 0: 	 branch_block_stmt_28/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/branch_block_stmt_28__entry__
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80__entry__
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_complete/req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_update_start_
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_update_start_
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_complete/req
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_update_start_
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/word_access_complete/word_0/cr
      -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_51_load_0_req_0); -- 
    cr_58_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_58_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_51_load_0_req_1); -- 
    req_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_74_index_offset_req_0); -- 
    req_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_60_index_offset_req_0); -- 
    req_94_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_94_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_60_index_offset_req_1); -- 
    req_109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_61_final_reg_req_1); -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_65_load_0_req_1); -- 
    req_190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_74_index_offset_req_1); -- 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_75_final_reg_req_1); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_79_load_0_req_1); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	316 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_28/$exit
      -- CP-element group 1: 	 branch_block_stmt_28/branch_block_stmt_28__exit__
      -- CP-element group 1: 	 branch_block_stmt_28/do_while_stmt_81__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(316);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/word_access_start/$exit
      -- CP-element group 2: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/word_access_start/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Sample/word_access_start/word_0/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_51_load_0_ack_0, ack => access_T_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	16 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/word_access_complete/$exit
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/word_access_complete/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/word_access_complete/word_0/ca
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/ptr_deref_51_Merge/$entry
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/ptr_deref_51_Merge/$exit
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/ptr_deref_51_Merge/merge_req
      -- CP-element group 3: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_51_Update/ptr_deref_51_Merge/merge_ack
      -- 
    ca_59_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_51_load_0_ack_1, ack => access_T_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	16 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_sample_complete
      -- CP-element group 4: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Sample/ack
      -- 
    ack_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_60_index_offset_ack_0, ack => access_T_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (11) 
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_root_address_calculated
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_offset_calculated
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_final_index_sum_regn_Update/ack
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_base_plus_offset/$entry
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_base_plus_offset/$exit
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_base_plus_offset/sum_rename_req
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_60_base_plus_offset/sum_rename_ack
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_request/$entry
      -- CP-element group 5: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_request/req
      -- 
    ack_95_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_60_index_offset_ack_1, ack => access_T_CP_0_elements(5)); -- 
    req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(5), ack => addr_of_61_final_reg_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_request/$exit
      -- CP-element group 6: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_request/ack
      -- 
    ack_105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_61_final_reg_ack_0, ack => access_T_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (24) 
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_61_complete/ack
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_word_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_root_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_address_resized
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_addr_resize/$entry
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_addr_resize/$exit
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_addr_resize/base_resize_req
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_addr_resize/base_resize_ack
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_plus_offset/$entry
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_plus_offset/$exit
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_plus_offset/sum_rename_req
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_base_plus_offset/sum_rename_ack
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_word_addrgen/$entry
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_word_addrgen/$exit
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_word_addrgen/root_register_req
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_word_addrgen/root_register_ack
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/word_access_start/word_0/rr
      -- 
    ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_61_final_reg_ack_1, ack => access_T_CP_0_elements(7)); -- 
    rr_143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(7), ack => ptr_deref_65_load_0_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/word_access_start/$exit
      -- CP-element group 8: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Sample/word_access_start/word_0/ra
      -- 
    ra_144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_65_load_0_ack_0, ack => access_T_CP_0_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/ptr_deref_65_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/ptr_deref_65_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/ptr_deref_65_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_65_Update/ptr_deref_65_Merge/merge_ack
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_65_load_0_ack_1, ack => access_T_CP_0_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	16 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_sample_complete
      -- CP-element group 10: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Sample/ack
      -- 
    ack_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_74_index_offset_ack_0, ack => access_T_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (11) 
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_offset_calculated
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_final_index_sum_regn_Update/ack
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_base_plus_offset/$entry
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_base_plus_offset/$exit
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_base_plus_offset/sum_rename_req
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/array_obj_ref_74_base_plus_offset/sum_rename_ack
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_request/$entry
      -- CP-element group 11: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_request/req
      -- 
    ack_191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_74_index_offset_ack_1, ack => access_T_CP_0_elements(11)); -- 
    req_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(11), ack => addr_of_75_final_reg_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_request/$exit
      -- CP-element group 12: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_request/ack
      -- 
    ack_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_75_final_reg_ack_0, ack => access_T_CP_0_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (24) 
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/addr_of_75_complete/ack
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_address_resized
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_addr_resize/$entry
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_addr_resize/$exit
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_addr_resize/base_resize_req
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_addr_resize/base_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_word_addrgen/root_register_ack
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/word_access_start/$entry
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/word_access_start/word_0/rr
      -- 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_75_final_reg_ack_1, ack => access_T_CP_0_elements(13)); -- 
    rr_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(13), ack => ptr_deref_79_load_0_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Sample/word_access_start/word_0/ra
      -- 
    ra_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_79_load_0_ack_0, ack => access_T_CP_0_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/ptr_deref_79_Merge/$entry
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/ptr_deref_79_Merge/$exit
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/ptr_deref_79_Merge/merge_req
      -- CP-element group 15: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/ptr_deref_79_Update/ptr_deref_79_Merge/merge_ack
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_79_load_0_ack_1, ack => access_T_CP_0_elements(15)); -- 
    -- CP-element group 16:  join  transition  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	4 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	10 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80/$exit
      -- CP-element group 16: 	 branch_block_stmt_28/assign_stmt_35_to_assign_stmt_80__exit__
      -- CP-element group 16: 	 branch_block_stmt_28/do_while_stmt_81__entry__
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(3) & access_T_CP_0_elements(4) & access_T_CP_0_elements(9) & access_T_CP_0_elements(10) & access_T_CP_0_elements(15);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	23 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_28/do_while_stmt_81/$entry
      -- CP-element group 17: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81__entry__
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(16);
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	316 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81__exit__
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  merge  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_28/do_while_stmt_81/loop_back
      -- 
    -- Element group access_T_CP_0_elements(19) is bound as output of CP function.
    -- CP-element group 20:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	25 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	314 
    -- CP-element group 20: 	315 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_81/condition_done
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_81/loop_exit/$entry
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_81/loop_taken/$entry
      -- 
    access_T_CP_0_elements(20) <= access_T_CP_0_elements(25);
    -- CP-element group 21:  branch  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	313 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_28/do_while_stmt_81/loop_body_done
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(313);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	133 
    -- CP-element group 22: 	116 
    -- CP-element group 22: 	97 
    -- CP-element group 22: 	36 
    -- CP-element group 22: 	55 
    -- CP-element group 22: 	76 
    -- CP-element group 22: 	152 
    -- CP-element group 22: 	171 
    -- CP-element group 22: 	190 
    -- CP-element group 22: 	209 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(22) <= access_T_CP_0_elements(19);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	135 
    -- CP-element group 23: 	118 
    -- CP-element group 23: 	99 
    -- CP-element group 23: 	38 
    -- CP-element group 23: 	57 
    -- CP-element group 23: 	78 
    -- CP-element group 23: 	154 
    -- CP-element group 23: 	173 
    -- CP-element group 23: 	192 
    -- CP-element group 23: 	211 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(17);
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	129 
    -- CP-element group 24: 	130 
    -- CP-element group 24: 	110 
    -- CP-element group 24: 	92 
    -- CP-element group 24: 	111 
    -- CP-element group 24: 	91 
    -- CP-element group 24: 	30 
    -- CP-element group 24: 	31 
    -- CP-element group 24: 	49 
    -- CP-element group 24: 	50 
    -- CP-element group 24: 	70 
    -- CP-element group 24: 	71 
    -- CP-element group 24: 	146 
    -- CP-element group 24: 	147 
    -- CP-element group 24: 	165 
    -- CP-element group 24: 	166 
    -- CP-element group 24: 	184 
    -- CP-element group 24: 	185 
    -- CP-element group 24: 	203 
    -- CP-element group 24: 	204 
    -- CP-element group 24: 	227 
    -- CP-element group 24: 	228 
    -- CP-element group 24: 	257 
    -- CP-element group 24: 	258 
    -- CP-element group 24: 	287 
    -- CP-element group 24: 	288 
    -- CP-element group 24: 	312 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/$entry
      -- CP-element group 24: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	96 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	170 
    -- CP-element group 25: 	312 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	20 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/condition_evaluated
      -- 
    condition_evaluated_271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(25), ack => do_while_stmt_81_branch_req_0); -- 
    access_T_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(96) & access_T_CP_0_elements(29) & access_T_CP_0_elements(170) & access_T_CP_0_elements(312);
      gj_access_T_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	129 
    -- CP-element group 26: 	110 
    -- CP-element group 26: 	91 
    -- CP-element group 26: 	30 
    -- CP-element group 26: 	49 
    -- CP-element group 26: 	70 
    -- CP-element group 26: 	146 
    -- CP-element group 26: 	165 
    -- CP-element group 26: 	184 
    -- CP-element group 26: 	203 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	29 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	93 
    -- CP-element group 26: 	112 
    -- CP-element group 26: 	32 
    -- CP-element group 26: 	51 
    -- CP-element group 26: 	72 
    -- CP-element group 26: 	148 
    -- CP-element group 26: 	167 
    -- CP-element group 26: 	186 
    -- CP-element group 26: 	205 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/aggregated_phi_sample_req
      -- CP-element group 26: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_sample_start__ps
      -- 
    access_T_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(129) & access_T_CP_0_elements(110) & access_T_CP_0_elements(91) & access_T_CP_0_elements(30) & access_T_CP_0_elements(49) & access_T_CP_0_elements(70) & access_T_CP_0_elements(146) & access_T_CP_0_elements(165) & access_T_CP_0_elements(184) & access_T_CP_0_elements(203) & access_T_CP_0_elements(29);
      gj_access_T_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	131 
    -- CP-element group 27: 	94 
    -- CP-element group 27: 	113 
    -- CP-element group 27: 	33 
    -- CP-element group 27: 	52 
    -- CP-element group 27: 	73 
    -- CP-element group 27: 	149 
    -- CP-element group 27: 	168 
    -- CP-element group 27: 	187 
    -- CP-element group 27: 	206 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	238 
    -- CP-element group 27: 	242 
    -- CP-element group 27: 	246 
    -- CP-element group 27: 	268 
    -- CP-element group 27: 	272 
    -- CP-element group 27: 	276 
    -- CP-element group 27: 	298 
    -- CP-element group 27: 	302 
    -- CP-element group 27: 	306 
    -- CP-element group 27: 	313 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	129 
    -- CP-element group 27: 	110 
    -- CP-element group 27: 	91 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	49 
    -- CP-element group 27: 	70 
    -- CP-element group 27: 	146 
    -- CP-element group 27: 	165 
    -- CP-element group 27: 	184 
    -- CP-element group 27: 	203 
    -- CP-element group 27:  members (11) 
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/aggregated_phi_sample_ack
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_sample_completed_
      -- 
    access_T_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= access_T_CP_0_elements(131) & access_T_CP_0_elements(94) & access_T_CP_0_elements(113) & access_T_CP_0_elements(33) & access_T_CP_0_elements(52) & access_T_CP_0_elements(73) & access_T_CP_0_elements(149) & access_T_CP_0_elements(168) & access_T_CP_0_elements(187) & access_T_CP_0_elements(206);
      gj_access_T_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	130 
    -- CP-element group 28: 	92 
    -- CP-element group 28: 	111 
    -- CP-element group 28: 	31 
    -- CP-element group 28: 	50 
    -- CP-element group 28: 	71 
    -- CP-element group 28: 	147 
    -- CP-element group 28: 	166 
    -- CP-element group 28: 	185 
    -- CP-element group 28: 	204 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	95 
    -- CP-element group 28: 	114 
    -- CP-element group 28: 	34 
    -- CP-element group 28: 	53 
    -- CP-element group 28: 	74 
    -- CP-element group 28: 	150 
    -- CP-element group 28: 	169 
    -- CP-element group 28: 	188 
    -- CP-element group 28: 	207 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/aggregated_phi_update_req
      -- CP-element group 28: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_update_start__ps
      -- 
    access_T_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= access_T_CP_0_elements(130) & access_T_CP_0_elements(92) & access_T_CP_0_elements(111) & access_T_CP_0_elements(31) & access_T_CP_0_elements(50) & access_T_CP_0_elements(71) & access_T_CP_0_elements(147) & access_T_CP_0_elements(166) & access_T_CP_0_elements(185) & access_T_CP_0_elements(204);
      gj_access_T_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	132 
    -- CP-element group 29: 	96 
    -- CP-element group 29: 	115 
    -- CP-element group 29: 	35 
    -- CP-element group 29: 	54 
    -- CP-element group 29: 	75 
    -- CP-element group 29: 	151 
    -- CP-element group 29: 	170 
    -- CP-element group 29: 	189 
    -- CP-element group 29: 	208 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	26 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= access_T_CP_0_elements(132) & access_T_CP_0_elements(96) & access_T_CP_0_elements(115) & access_T_CP_0_elements(35) & access_T_CP_0_elements(54) & access_T_CP_0_elements(75) & access_T_CP_0_elements(151) & access_T_CP_0_elements(170) & access_T_CP_0_elements(189) & access_T_CP_0_elements(208);
      gj_access_T_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	26 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_sample_start_
      -- 
    access_T_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	24 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	35 
    -- CP-element group 31: 	229 
    -- CP-element group 31: 	235 
    -- CP-element group 31: 	243 
    -- CP-element group 31: 	250 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	28 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_update_start_
      -- 
    access_T_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(35) & access_T_CP_0_elements(229) & access_T_CP_0_elements(235) & access_T_CP_0_elements(243) & access_T_CP_0_elements(250);
      gj_access_T_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	26 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_sample_start__ps
      -- 
    access_T_CP_0_elements(32) <= access_T_CP_0_elements(26);
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	27 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(33) is bound as output of CP function.
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	28 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_update_start__ps
      -- 
    access_T_CP_0_elements(34) <= access_T_CP_0_elements(28);
    -- CP-element group 35:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	29 
    -- CP-element group 35: 	229 
    -- CP-element group 35: 	233 
    -- CP-element group 35: 	241 
    -- CP-element group 35: 	249 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	31 
    -- CP-element group 35:  members (15) 
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Sample/req
      -- 
    req_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(35), ack => array_obj_ref_197_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	22 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_loopback_trigger
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(22);
    -- CP-element group 37:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_loopback_sample_req
      -- CP-element group 37: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_loopback_sample_req_ps
      -- 
    phi_stmt_83_loopback_sample_req_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_83_loopback_sample_req_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(37), ack => phi_stmt_83_req_1); -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	23 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_entry_trigger
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(23);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_entry_sample_req
      -- CP-element group 39: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_entry_sample_req_ps
      -- 
    phi_stmt_83_entry_sample_req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_83_entry_sample_req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(39), ack => phi_stmt_83_req_0); -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_phi_mux_ack
      -- CP-element group 40: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_83_phi_mux_ack_ps
      -- 
    phi_stmt_83_phi_mux_ack_292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_83_ack_0, ack => access_T_CP_0_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_sample_start__ps
      -- CP-element group 41: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_sample_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_update_start__ps
      -- CP-element group 42: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_update_start_
      -- 
    -- Element group access_T_CP_0_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_update_completed__ps
      -- 
    access_T_CP_0_elements(43) <= access_T_CP_0_elements(44);
    -- CP-element group 44:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	43 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_86_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(44) is a control-delay.
    cp_element_44_delay: control_delay_element  generic map(name => " 44_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(42), ack => access_T_CP_0_elements(44), clk => clk, reset =>reset);
    -- CP-element group 45:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Sample/req
      -- 
    req_313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(45), ack => n_address1_176_87_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_update_start_
      -- CP-element group 46: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Update/req
      -- 
    req_318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(46), ack => n_address1_176_87_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Sample/ack
      -- 
    ack_314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_176_87_buf_ack_0, ack => access_T_CP_0_elements(47)); -- 
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_update_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address1_87_Update/ack
      -- 
    ack_319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_176_87_buf_ack_1, ack => access_T_CP_0_elements(48)); -- 
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	24 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	27 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	26 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_sample_start_
      -- 
    access_T_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	24 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	54 
    -- CP-element group 50: 	259 
    -- CP-element group 50: 	265 
    -- CP-element group 50: 	273 
    -- CP-element group 50: 	280 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	28 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_update_start_
      -- 
    access_T_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(54) & access_T_CP_0_elements(259) & access_T_CP_0_elements(265) & access_T_CP_0_elements(273) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	26 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_sample_start__ps
      -- 
    access_T_CP_0_elements(51) <= access_T_CP_0_elements(26);
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	27 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(52) is bound as output of CP function.
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	28 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_update_start__ps
      -- 
    access_T_CP_0_elements(53) <= access_T_CP_0_elements(28);
    -- CP-element group 54:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	29 
    -- CP-element group 54: 	259 
    -- CP-element group 54: 	263 
    -- CP-element group 54: 	271 
    -- CP-element group 54: 	279 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	50 
    -- CP-element group 54:  members (15) 
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_computed_1
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_scaled_1
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_resized_1
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Sample/req
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_scale_1/scale_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_scale_1/scale_rename_req
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_scale_1/$exit
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_scale_1/$entry
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_resize_1/index_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_resize_1/index_resize_req
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_resize_1/$exit
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_index_resize_1/$entry
      -- 
    req_971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(54), ack => array_obj_ref_271_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	22 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_loopback_trigger
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(22);
    -- CP-element group 56:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_loopback_sample_req
      -- CP-element group 56: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_loopback_sample_req_ps
      -- 
    phi_stmt_88_loopback_sample_req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_88_loopback_sample_req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(56), ack => phi_stmt_88_req_1); -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	23 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_entry_trigger
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(23);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_entry_sample_req
      -- CP-element group 58: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_entry_sample_req_ps
      -- 
    phi_stmt_88_entry_sample_req_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_88_entry_sample_req_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(58), ack => phi_stmt_88_req_0); -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_phi_mux_ack
      -- CP-element group 59: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_88_phi_mux_ack_ps
      -- 
    phi_stmt_88_phi_mux_ack_336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_88_ack_0, ack => access_T_CP_0_elements(59)); -- 
    -- CP-element group 60:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Sample/rr
      -- 
    rr_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => type_cast_91_inst_req_0); -- 
    access_T_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(60) & access_T_CP_0_elements(64);
      gj_access_T_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_update_start_
      -- CP-element group 63: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Update/cr
      -- 
    cr_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(63), ack => type_cast_91_inst_req_1); -- 
    access_T_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(61) & access_T_CP_0_elements(65);
      gj_access_T_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Sample/ra
      -- 
    ra_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_91_inst_ack_0, ack => access_T_CP_0_elements(64)); -- 
    -- CP-element group 65:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_update_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_91_Update/ca
      -- 
    ca_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_91_inst_ack_1, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Sample/req
      -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(66), ack => n_address2_250_92_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_update_start_
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Update/req
      -- 
    req_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(67), ack => n_address2_250_92_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Sample/ack
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_250_92_buf_ack_0, ack => access_T_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address2_92_Update/ack
      -- 
    ack_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_250_92_buf_ack_1, ack => access_T_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	24 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	27 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	26 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_sample_start_
      -- 
    access_T_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	24 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	75 
    -- CP-element group 71: 	289 
    -- CP-element group 71: 	295 
    -- CP-element group 71: 	303 
    -- CP-element group 71: 	310 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	28 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_update_start_
      -- 
    access_T_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(75) & access_T_CP_0_elements(289) & access_T_CP_0_elements(295) & access_T_CP_0_elements(303) & access_T_CP_0_elements(310);
      gj_access_T_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	26 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_sample_start__ps
      -- 
    access_T_CP_0_elements(72) <= access_T_CP_0_elements(26);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	27 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_update_start__ps
      -- 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(28);
    -- CP-element group 75:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	29 
    -- CP-element group 75: 	289 
    -- CP-element group 75: 	293 
    -- CP-element group 75: 	301 
    -- CP-element group 75: 	309 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	71 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_scale_1/scale_rename_req
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_scale_1/scale_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_scale_1/$exit
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_scale_1/$entry
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_resize_1/index_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_resize_1/index_resize_req
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_resize_1/$exit
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_resize_1/$entry
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_computed_1
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_scaled_1
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_index_resized_1
      -- 
    req_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(75), ack => array_obj_ref_350_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	22 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_loopback_trigger
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(22);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_loopback_sample_req_ps
      -- 
    phi_stmt_93_loopback_sample_req_384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_93_loopback_sample_req_384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(77), ack => phi_stmt_93_req_1); -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	23 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_entry_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(23);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_entry_sample_req_ps
      -- 
    phi_stmt_93_entry_sample_req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_93_entry_sample_req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_93_req_0); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_93_phi_mux_ack_ps
      -- 
    phi_stmt_93_phi_mux_ack_390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_93_ack_0, ack => access_T_CP_0_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Sample/rr
      -- 
    rr_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => type_cast_96_inst_req_0); -- 
    access_T_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(85);
      gj_access_T_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_update_start_
      -- CP-element group 84: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Update/cr
      -- 
    cr_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(84), ack => type_cast_96_inst_req_1); -- 
    access_T_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(82) & access_T_CP_0_elements(86);
      gj_access_T_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Sample/ra
      -- 
    ra_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_0, ack => access_T_CP_0_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_96_Update/ca
      -- 
    ca_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_1, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Sample/req
      -- 
    req_421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(87), ack => n_address3_324_97_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_update_start_
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Update/req
      -- 
    req_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => n_address3_324_97_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Sample/ack
      -- 
    ack_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_324_97_buf_ack_0, ack => access_T_CP_0_elements(89)); -- 
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_address3_97_Update/ack
      -- 
    ack_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_324_97_buf_ack_1, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	24 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	27 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	26 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_sample_start_
      -- 
    access_T_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	24 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	96 
    -- CP-element group 92: 	224 
    -- CP-element group 92: 	254 
    -- CP-element group 92: 	284 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	28 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_update_start_
      -- 
    access_T_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(96) & access_T_CP_0_elements(224) & access_T_CP_0_elements(254) & access_T_CP_0_elements(284);
      gj_access_T_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	26 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_sample_start__ps
      -- 
    access_T_CP_0_elements(93) <= access_T_CP_0_elements(26);
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	27 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	28 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_update_start__ps
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(28);
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	25 
    -- CP-element group 96: 	29 
    -- CP-element group 96: 	222 
    -- CP-element group 96: 	252 
    -- CP-element group 96: 	282 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	92 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	22 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_loopback_trigger
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(22);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_loopback_sample_req
      -- CP-element group 98: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_loopback_sample_req_ps
      -- 
    phi_stmt_98_loopback_sample_req_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_98_loopback_sample_req_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => phi_stmt_98_req_1); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	23 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_entry_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(23);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_entry_sample_req
      -- CP-element group 100: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_entry_sample_req_ps
      -- 
    phi_stmt_98_entry_sample_req_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_98_entry_sample_req_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_98_req_0); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_phi_mux_ack
      -- CP-element group 101: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_98_phi_mux_ack_ps
      -- 
    phi_stmt_98_phi_mux_ack_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_98_ack_0, ack => access_T_CP_0_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_sample_start__ps
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_sample_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_update_start__ps
      -- CP-element group 103: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_update_start_
      -- 
    -- Element group access_T_CP_0_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_update_completed__ps
      -- 
    access_T_CP_0_elements(104) <= access_T_CP_0_elements(105);
    -- CP-element group 105:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	104 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_101_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(103), ack => access_T_CP_0_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Sample/req
      -- 
    req_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(106), ack => n_mycounter_143_102_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_update_start_
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Update/req
      -- 
    req_470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(107), ack => n_mycounter_143_102_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Sample/ack
      -- 
    ack_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_143_102_buf_ack_0, ack => access_T_CP_0_elements(108)); -- 
    -- CP-element group 109:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_update_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_mycounter_102_Update/ack
      -- 
    ack_471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_143_102_buf_ack_1, ack => access_T_CP_0_elements(109)); -- 
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	24 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	27 
    -- CP-element group 110: 	240 
    -- CP-element group 110: 	244 
    -- CP-element group 110: 	248 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	26 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_sample_start_
      -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27) & access_T_CP_0_elements(240) & access_T_CP_0_elements(244) & access_T_CP_0_elements(248);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	24 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	115 
    -- CP-element group 111: 	247 
    -- CP-element group 111: 	250 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	28 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_update_start_
      -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(115) & access_T_CP_0_elements(247) & access_T_CP_0_elements(250);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	26 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_sample_start__ps
      -- 
    access_T_CP_0_elements(112) <= access_T_CP_0_elements(26);
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	27 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	28 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_update_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(28);
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	29 
    -- CP-element group 115: 	245 
    -- CP-element group 115: 	249 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	111 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	22 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_loopback_trigger
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(22);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_loopback_sample_req
      -- CP-element group 117: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_loopback_sample_req_ps
      -- 
    phi_stmt_103_loopback_sample_req_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_103_loopback_sample_req_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_103_req_1); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	23 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_entry_trigger
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(23);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_entry_sample_req
      -- CP-element group 119: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_entry_sample_req_ps
      -- 
    phi_stmt_103_entry_sample_req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_103_entry_sample_req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_103_req_0); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_phi_mux_ack
      -- CP-element group 120: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_103_phi_mux_ack_ps
      -- 
    phi_stmt_103_phi_mux_ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_103_ack_0, ack => access_T_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Sample/req
      -- 
    req_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(121), ack => my_fetch1_52_105_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_update_start_
      -- CP-element group 122: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Update/req
      -- 
    req_506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(122), ack => my_fetch1_52_105_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_sample_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Sample/ack
      -- 
    ack_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_52_105_buf_ack_0, ack => access_T_CP_0_elements(123)); -- 
    -- CP-element group 124:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_update_completed__ps
      -- CP-element group 124: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch1_105_Update/ack
      -- 
    ack_507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_52_105_buf_ack_1, ack => access_T_CP_0_elements(124)); -- 
    -- CP-element group 125:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Sample/req
      -- 
    req_519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => n_fetch_val1_219_106_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_update_start_
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Update/req
      -- 
    req_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(126), ack => n_fetch_val1_219_106_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Sample/ack
      -- 
    ack_520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_219_106_buf_ack_0, ack => access_T_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_update_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val1_106_Update/ack
      -- 
    ack_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_219_106_buf_ack_1, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	24 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	27 
    -- CP-element group 129: 	270 
    -- CP-element group 129: 	274 
    -- CP-element group 129: 	278 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	26 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_sample_start_
      -- 
    access_T_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27) & access_T_CP_0_elements(270) & access_T_CP_0_elements(274) & access_T_CP_0_elements(278);
      gj_access_T_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	24 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: 	277 
    -- CP-element group 130: 	280 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	28 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_update_start_
      -- 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(132) & access_T_CP_0_elements(277) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	27 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(131) is bound as output of CP function.
    -- CP-element group 132:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	29 
    -- CP-element group 132: 	275 
    -- CP-element group 132: 	279 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	130 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	22 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_loopback_trigger
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(22);
    -- CP-element group 134:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_loopback_sample_req
      -- CP-element group 134: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_loopback_sample_req_ps
      -- 
    phi_stmt_107_loopback_sample_req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_loopback_sample_req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(134), ack => phi_stmt_107_req_1); -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	23 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_entry_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(23);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_entry_sample_req
      -- CP-element group 136: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_entry_sample_req_ps
      -- 
    phi_stmt_107_entry_sample_req_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_entry_sample_req_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_107_req_0); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (2) 
      -- CP-element group 137: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_phi_mux_ack
      -- CP-element group 137: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_107_phi_mux_ack_ps
      -- 
    phi_stmt_107_phi_mux_ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_107_ack_0, ack => access_T_CP_0_elements(137)); -- 
    -- CP-element group 138:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_sample_start__ps
      -- CP-element group 138: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Sample/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => my_fetch2_66_109_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_update_start__ps
      -- CP-element group 139: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_update_start_
      -- CP-element group 139: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Update/req
      -- 
    req_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(139), ack => my_fetch2_66_109_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(139) is bound as output of CP function.
    -- CP-element group 140:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Sample/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_66_109_buf_ack_0, ack => access_T_CP_0_elements(140)); -- 
    -- CP-element group 141:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_update_completed__ps
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch2_109_Update/ack
      -- 
    ack_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_66_109_buf_ack_1, ack => access_T_CP_0_elements(141)); -- 
    -- CP-element group 142:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_sample_start__ps
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Sample/req
      -- 
    req_573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(142), ack => n_fetch_val2_293_110_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(142) is bound as output of CP function.
    -- CP-element group 143:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_update_start__ps
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_update_start_
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Update/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(143), ack => n_fetch_val2_293_110_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(143) is bound as output of CP function.
    -- CP-element group 144:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_sample_completed__ps
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Sample/ack
      -- 
    ack_574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_293_110_buf_ack_0, ack => access_T_CP_0_elements(144)); -- 
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (4) 
      -- CP-element group 145: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_update_completed__ps
      -- CP-element group 145: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val2_110_Update/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_293_110_buf_ack_1, ack => access_T_CP_0_elements(145)); -- 
    -- CP-element group 146:  join  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	24 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	27 
    -- CP-element group 146: 	300 
    -- CP-element group 146: 	304 
    -- CP-element group 146: 	308 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	26 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_sample_start_
      -- 
    access_T_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	24 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	151 
    -- CP-element group 147: 	307 
    -- CP-element group 147: 	310 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	28 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_update_start_
      -- 
    access_T_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(151) & access_T_CP_0_elements(307) & access_T_CP_0_elements(310);
      gj_access_T_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	26 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_sample_start__ps
      -- 
    access_T_CP_0_elements(148) <= access_T_CP_0_elements(26);
    -- CP-element group 149:  join  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	27 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(149) is bound as output of CP function.
    -- CP-element group 150:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	28 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_update_start__ps
      -- 
    access_T_CP_0_elements(150) <= access_T_CP_0_elements(28);
    -- CP-element group 151:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	29 
    -- CP-element group 151: 	305 
    -- CP-element group 151: 	309 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	147 
    -- CP-element group 151:  members (2) 
      -- CP-element group 151: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(151) is bound as output of CP function.
    -- CP-element group 152:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	22 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (1) 
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_loopback_trigger
      -- 
    access_T_CP_0_elements(152) <= access_T_CP_0_elements(22);
    -- CP-element group 153:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_loopback_sample_req
      -- CP-element group 153: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_loopback_sample_req_ps
      -- 
    phi_stmt_111_loopback_sample_req_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_111_loopback_sample_req_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(153), ack => phi_stmt_111_req_1); -- 
    -- Element group access_T_CP_0_elements(153) is bound as output of CP function.
    -- CP-element group 154:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	23 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_entry_trigger
      -- 
    access_T_CP_0_elements(154) <= access_T_CP_0_elements(23);
    -- CP-element group 155:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (2) 
      -- CP-element group 155: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_entry_sample_req
      -- CP-element group 155: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_entry_sample_req_ps
      -- 
    phi_stmt_111_entry_sample_req_593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_111_entry_sample_req_593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => phi_stmt_111_req_0); -- 
    -- Element group access_T_CP_0_elements(155) is bound as output of CP function.
    -- CP-element group 156:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_phi_mux_ack
      -- CP-element group 156: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_111_phi_mux_ack_ps
      -- 
    phi_stmt_111_phi_mux_ack_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_111_ack_0, ack => access_T_CP_0_elements(156)); -- 
    -- CP-element group 157:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (4) 
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_sample_start__ps
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Sample/req
      -- 
    req_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(157), ack => my_fetch3_80_113_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(157) is bound as output of CP function.
    -- CP-element group 158:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (4) 
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_update_start__ps
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_update_start_
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Update/req
      -- 
    req_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(158), ack => my_fetch3_80_113_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(158) is bound as output of CP function.
    -- CP-element group 159:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (4) 
      -- CP-element group 159: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_sample_completed__ps
      -- CP-element group 159: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Sample/ack
      -- 
    ack_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_80_113_buf_ack_0, ack => access_T_CP_0_elements(159)); -- 
    -- CP-element group 160:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (4) 
      -- CP-element group 160: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_update_completed__ps
      -- CP-element group 160: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_my_fetch3_113_Update/ack
      -- 
    ack_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_80_113_buf_ack_1, ack => access_T_CP_0_elements(160)); -- 
    -- CP-element group 161:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (4) 
      -- CP-element group 161: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_sample_start__ps
      -- CP-element group 161: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Sample/req
      -- 
    req_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(161), ack => n_fetch_val3_372_114_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(161) is bound as output of CP function.
    -- CP-element group 162:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (4) 
      -- CP-element group 162: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_update_start__ps
      -- CP-element group 162: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_update_start_
      -- CP-element group 162: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Update/req
      -- 
    req_632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(162), ack => n_fetch_val3_372_114_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(162) is bound as output of CP function.
    -- CP-element group 163:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (4) 
      -- CP-element group 163: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_sample_completed__ps
      -- CP-element group 163: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Sample/ack
      -- 
    ack_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_372_114_buf_ack_0, ack => access_T_CP_0_elements(163)); -- 
    -- CP-element group 164:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (4) 
      -- CP-element group 164: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_update_completed__ps
      -- CP-element group 164: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_fetch_val3_114_Update/ack
      -- 
    ack_633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_372_114_buf_ack_1, ack => access_T_CP_0_elements(164)); -- 
    -- CP-element group 165:  join  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	24 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	27 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	26 
    -- CP-element group 165:  members (1) 
      -- CP-element group 165: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_sample_start_
      -- 
    access_T_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	24 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	170 
    -- CP-element group 166: 	224 
    -- CP-element group 166: 	254 
    -- CP-element group 166: 	284 
    -- CP-element group 166: 	310 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	28 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_update_start_
      -- 
    access_T_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(170) & access_T_CP_0_elements(224) & access_T_CP_0_elements(254) & access_T_CP_0_elements(284) & access_T_CP_0_elements(310);
      gj_access_T_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	26 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_sample_start__ps
      -- 
    access_T_CP_0_elements(167) <= access_T_CP_0_elements(26);
    -- CP-element group 168:  join  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	27 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(168) is bound as output of CP function.
    -- CP-element group 169:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	28 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (1) 
      -- CP-element group 169: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_update_start__ps
      -- 
    access_T_CP_0_elements(169) <= access_T_CP_0_elements(28);
    -- CP-element group 170:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	25 
    -- CP-element group 170: 	29 
    -- CP-element group 170: 	222 
    -- CP-element group 170: 	252 
    -- CP-element group 170: 	282 
    -- CP-element group 170: 	309 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	166 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(170) is bound as output of CP function.
    -- CP-element group 171:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	22 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_loopback_trigger
      -- 
    access_T_CP_0_elements(171) <= access_T_CP_0_elements(22);
    -- CP-element group 172:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_loopback_sample_req
      -- CP-element group 172: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_loopback_sample_req_ps
      -- 
    phi_stmt_115_loopback_sample_req_644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_115_loopback_sample_req_644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => phi_stmt_115_req_1); -- 
    -- Element group access_T_CP_0_elements(172) is bound as output of CP function.
    -- CP-element group 173:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	23 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_entry_trigger
      -- 
    access_T_CP_0_elements(173) <= access_T_CP_0_elements(23);
    -- CP-element group 174:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (2) 
      -- CP-element group 174: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_entry_sample_req
      -- CP-element group 174: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_entry_sample_req_ps
      -- 
    phi_stmt_115_entry_sample_req_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_115_entry_sample_req_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(174), ack => phi_stmt_115_req_0); -- 
    -- Element group access_T_CP_0_elements(174) is bound as output of CP function.
    -- CP-element group 175:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (2) 
      -- CP-element group 175: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_phi_mux_ack
      -- CP-element group 175: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_115_phi_mux_ack_ps
      -- 
    phi_stmt_115_phi_mux_ack_650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_115_ack_0, ack => access_T_CP_0_elements(175)); -- 
    -- CP-element group 176:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (4) 
      -- CP-element group 176: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_sample_start__ps
      -- CP-element group 176: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_sample_completed__ps
      -- CP-element group 176: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(176) is bound as output of CP function.
    -- CP-element group 177:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (2) 
      -- CP-element group 177: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_update_start__ps
      -- CP-element group 177: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_update_start_
      -- 
    -- Element group access_T_CP_0_elements(177) is bound as output of CP function.
    -- CP-element group 178:  join  transition  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (1) 
      -- CP-element group 178: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_update_completed__ps
      -- 
    access_T_CP_0_elements(178) <= access_T_CP_0_elements(179);
    -- CP-element group 179:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	178 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_118_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(179) is a control-delay.
    cp_element_179_delay: control_delay_element  generic map(name => " 179_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(177), ack => access_T_CP_0_elements(179), clk => clk, reset =>reset);
    -- CP-element group 180:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (4) 
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_sample_start__ps
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Sample/req
      -- 
    req_671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => n_row1_171_119_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(180) is bound as output of CP function.
    -- CP-element group 181:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (4) 
      -- CP-element group 181: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_update_start__ps
      -- CP-element group 181: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_update_start_
      -- CP-element group 181: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Update/req
      -- 
    req_676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(181), ack => n_row1_171_119_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(181) is bound as output of CP function.
    -- CP-element group 182:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (4) 
      -- CP-element group 182: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_sample_completed__ps
      -- CP-element group 182: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Sample/ack
      -- 
    ack_672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_171_119_buf_ack_0, ack => access_T_CP_0_elements(182)); -- 
    -- CP-element group 183:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (4) 
      -- CP-element group 183: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_update_completed__ps
      -- CP-element group 183: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row1_119_Update/ack
      -- 
    ack_677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_171_119_buf_ack_1, ack => access_T_CP_0_elements(183)); -- 
    -- CP-element group 184:  join  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	24 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	27 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	26 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_sample_start_
      -- 
    access_T_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	24 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	189 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	28 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_update_start_
      -- 
    access_T_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(189);
      gj_access_T_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	26 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_sample_start__ps
      -- 
    access_T_CP_0_elements(186) <= access_T_CP_0_elements(26);
    -- CP-element group 187:  join  transition  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	27 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(187) is bound as output of CP function.
    -- CP-element group 188:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	28 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_update_start__ps
      -- 
    access_T_CP_0_elements(188) <= access_T_CP_0_elements(28);
    -- CP-element group 189:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	29 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	185 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(189) is bound as output of CP function.
    -- CP-element group 190:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	22 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (1) 
      -- CP-element group 190: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_loopback_trigger
      -- 
    access_T_CP_0_elements(190) <= access_T_CP_0_elements(22);
    -- CP-element group 191:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (2) 
      -- CP-element group 191: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_loopback_sample_req
      -- CP-element group 191: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_loopback_sample_req_ps
      -- 
    phi_stmt_120_loopback_sample_req_688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_120_loopback_sample_req_688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(191), ack => phi_stmt_120_req_1); -- 
    -- Element group access_T_CP_0_elements(191) is bound as output of CP function.
    -- CP-element group 192:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	23 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_entry_trigger
      -- 
    access_T_CP_0_elements(192) <= access_T_CP_0_elements(23);
    -- CP-element group 193:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (2) 
      -- CP-element group 193: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_entry_sample_req
      -- CP-element group 193: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_entry_sample_req_ps
      -- 
    phi_stmt_120_entry_sample_req_691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_120_entry_sample_req_691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => phi_stmt_120_req_0); -- 
    -- Element group access_T_CP_0_elements(193) is bound as output of CP function.
    -- CP-element group 194:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (2) 
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_phi_mux_ack
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_120_phi_mux_ack_ps
      -- 
    phi_stmt_120_phi_mux_ack_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_120_ack_0, ack => access_T_CP_0_elements(194)); -- 
    -- CP-element group 195:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (4) 
      -- CP-element group 195: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_sample_start__ps
      -- CP-element group 195: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_sample_completed__ps
      -- CP-element group 195: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(195) is bound as output of CP function.
    -- CP-element group 196:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (2) 
      -- CP-element group 196: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_update_start__ps
      -- CP-element group 196: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_update_start_
      -- 
    -- Element group access_T_CP_0_elements(196) is bound as output of CP function.
    -- CP-element group 197:  join  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	198 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_update_completed__ps
      -- 
    access_T_CP_0_elements(197) <= access_T_CP_0_elements(198);
    -- CP-element group 198:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	197 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_123_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(198) is a control-delay.
    cp_element_198_delay: control_delay_element  generic map(name => " 198_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(196), ack => access_T_CP_0_elements(198), clk => clk, reset =>reset);
    -- CP-element group 199:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (4) 
      -- CP-element group 199: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_sample_start__ps
      -- CP-element group 199: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Sample/req
      -- 
    req_715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(199), ack => n_row2_245_124_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(199) is bound as output of CP function.
    -- CP-element group 200:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (4) 
      -- CP-element group 200: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_update_start__ps
      -- CP-element group 200: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_update_start_
      -- CP-element group 200: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Update/req
      -- 
    req_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => n_row2_245_124_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(200) is bound as output of CP function.
    -- CP-element group 201:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (4) 
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_sample_completed__ps
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Sample/ack
      -- 
    ack_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_245_124_buf_ack_0, ack => access_T_CP_0_elements(201)); -- 
    -- CP-element group 202:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (4) 
      -- CP-element group 202: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_update_completed__ps
      -- CP-element group 202: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row2_124_Update/ack
      -- 
    ack_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_245_124_buf_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  join  transition  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	24 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	27 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	26 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_sample_start_
      -- 
    access_T_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	24 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	208 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	28 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_update_start_
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(208);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	26 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_sample_start__ps
      -- 
    access_T_CP_0_elements(205) <= access_T_CP_0_elements(26);
    -- CP-element group 206:  join  transition  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	27 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(206) is bound as output of CP function.
    -- CP-element group 207:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	28 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_update_start__ps
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(28);
    -- CP-element group 208:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	29 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	204 
    -- CP-element group 208:  members (2) 
      -- CP-element group 208: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(208) is bound as output of CP function.
    -- CP-element group 209:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	22 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_loopback_trigger
      -- 
    access_T_CP_0_elements(209) <= access_T_CP_0_elements(22);
    -- CP-element group 210:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (2) 
      -- CP-element group 210: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_loopback_sample_req
      -- CP-element group 210: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_loopback_sample_req_ps
      -- 
    phi_stmt_125_loopback_sample_req_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_125_loopback_sample_req_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(210), ack => phi_stmt_125_req_1); -- 
    -- Element group access_T_CP_0_elements(210) is bound as output of CP function.
    -- CP-element group 211:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	23 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_entry_trigger
      -- 
    access_T_CP_0_elements(211) <= access_T_CP_0_elements(23);
    -- CP-element group 212:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (2) 
      -- CP-element group 212: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_entry_sample_req
      -- CP-element group 212: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_entry_sample_req_ps
      -- 
    phi_stmt_125_entry_sample_req_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_125_entry_sample_req_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(212), ack => phi_stmt_125_req_0); -- 
    -- Element group access_T_CP_0_elements(212) is bound as output of CP function.
    -- CP-element group 213:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (2) 
      -- CP-element group 213: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_phi_mux_ack
      -- CP-element group 213: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/phi_stmt_125_phi_mux_ack_ps
      -- 
    phi_stmt_125_phi_mux_ack_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_125_ack_0, ack => access_T_CP_0_elements(213)); -- 
    -- CP-element group 214:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (4) 
      -- CP-element group 214: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_sample_start__ps
      -- CP-element group 214: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_sample_completed__ps
      -- CP-element group 214: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(214) is bound as output of CP function.
    -- CP-element group 215:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (2) 
      -- CP-element group 215: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_update_start__ps
      -- CP-element group 215: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_update_start_
      -- 
    -- Element group access_T_CP_0_elements(215) is bound as output of CP function.
    -- CP-element group 216:  join  transition  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	217 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (1) 
      -- CP-element group 216: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_update_completed__ps
      -- 
    access_T_CP_0_elements(216) <= access_T_CP_0_elements(217);
    -- CP-element group 217:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	216 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/type_cast_128_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(217) is a control-delay.
    cp_element_217_delay: control_delay_element  generic map(name => " 217_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(215), ack => access_T_CP_0_elements(217), clk => clk, reset =>reset);
    -- CP-element group 218:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (4) 
      -- CP-element group 218: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_sample_start__ps
      -- CP-element group 218: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Sample/req
      -- 
    req_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(218), ack => n_row3_319_129_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(218) is bound as output of CP function.
    -- CP-element group 219:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (4) 
      -- CP-element group 219: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_update_start__ps
      -- CP-element group 219: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_update_start_
      -- CP-element group 219: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Update/req
      -- 
    req_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(219), ack => n_row3_319_129_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(219) is bound as output of CP function.
    -- CP-element group 220:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (4) 
      -- CP-element group 220: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_sample_completed__ps
      -- CP-element group 220: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Sample/ack
      -- 
    ack_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_319_129_buf_ack_0, ack => access_T_CP_0_elements(220)); -- 
    -- CP-element group 221:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (4) 
      -- CP-element group 221: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_update_completed__ps
      -- CP-element group 221: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/R_n_row3_129_Update/ack
      -- 
    ack_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_319_129_buf_ack_1, ack => access_T_CP_0_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	96 
    -- CP-element group 222: 	170 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Sample/req
      -- 
    req_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(222), ack => W_continue_185_delayed_1_0_177_inst_req_0); -- 
    access_T_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(96) & access_T_CP_0_elements(170) & access_T_CP_0_elements(224);
      gj_access_T_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	225 
    -- CP-element group 223: 	235 
    -- CP-element group 223: 	243 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_update_start_
      -- CP-element group 223: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Update/req
      -- 
    req_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(223), ack => W_continue_185_delayed_1_0_177_inst_req_1); -- 
    access_T_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(225) & access_T_CP_0_elements(235) & access_T_CP_0_elements(243);
      gj_access_T_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	92 
    -- CP-element group 224: 	166 
    -- CP-element group 224: 	222 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Sample/ack
      -- 
    ack_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_185_delayed_1_0_177_inst_ack_0, ack => access_T_CP_0_elements(224)); -- 
    -- CP-element group 225:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	233 
    -- CP-element group 225: 	241 
    -- CP-element group 225: marked-successors 
    -- CP-element group 225: 	223 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_179_Update/ack
      -- 
    ack_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_185_delayed_1_0_177_inst_ack_1, ack => access_T_CP_0_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	230 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	231 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	231 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_request/$entry
      -- CP-element group 226: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_request/req
      -- 
    req_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(226), ack => addr_of_198_final_reg_req_0); -- 
    access_T_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(230) & access_T_CP_0_elements(231);
      gj_access_T_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	24 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	232 
    -- CP-element group 227: 	239 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	232 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_update_start_
      -- CP-element group 227: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_complete/$entry
      -- CP-element group 227: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_complete/req
      -- 
    req_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(227), ack => addr_of_198_final_reg_req_1); -- 
    access_T_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(232) & access_T_CP_0_elements(239);
      gj_access_T_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	24 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: 	231 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_update_start
      -- CP-element group 228: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Update/req
      -- 
    req_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(228), ack => array_obj_ref_197_index_offset_req_1); -- 
    access_T_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(230) & access_T_CP_0_elements(231);
      gj_access_T_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	35 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	313 
    -- CP-element group 229: marked-successors 
    -- CP-element group 229: 	31 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_sample_complete
      -- CP-element group 229: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Sample/ack
      -- 
    ack_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_index_offset_ack_0, ack => access_T_CP_0_elements(229)); -- 
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	226 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (8) 
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_root_address_calculated
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_offset_calculated
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_final_index_sum_regn_Update/ack
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_base_plus_offset/$entry
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_base_plus_offset/$exit
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_base_plus_offset/sum_rename_req
      -- CP-element group 230: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_197_base_plus_offset/sum_rename_ack
      -- 
    ack_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_index_offset_ack_1, ack => access_T_CP_0_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	226 
    -- CP-element group 231: successors 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	226 
    -- CP-element group 231: 	228 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_request/$exit
      -- CP-element group 231: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_request/ack
      -- 
    ack_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_198_final_reg_ack_0, ack => access_T_CP_0_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	227 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	237 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	227 
    -- CP-element group 232:  members (19) 
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_complete/$exit
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_198_complete/ack
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_word_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_root_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_address_resized
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_addr_resize/$entry
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_addr_resize/$exit
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_addr_resize/base_resize_req
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_addr_resize/base_resize_ack
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_plus_offset/$entry
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_plus_offset/$exit
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_plus_offset/sum_rename_req
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_base_plus_offset/sum_rename_ack
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_word_addrgen/$entry
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_word_addrgen/$exit
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_word_addrgen/root_register_req
      -- CP-element group 232: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_word_addrgen/root_register_ack
      -- 
    ack_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_198_final_reg_ack_1, ack => access_T_CP_0_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	35 
    -- CP-element group 233: 	225 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Sample/req
      -- 
    req_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(233), ack => W_fn1_197_delayed_7_0_200_inst_req_0); -- 
    access_T_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(35) & access_T_CP_0_elements(225) & access_T_CP_0_elements(235);
      gj_access_T_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: 	239 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_update_start_
      -- CP-element group 234: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Update/req
      -- 
    req_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(234), ack => W_fn1_197_delayed_7_0_200_inst_req_1); -- 
    access_T_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(236) & access_T_CP_0_elements(239);
      gj_access_T_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	31 
    -- CP-element group 235: 	223 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Sample/ack
      -- 
    ack_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_197_delayed_7_0_200_inst_ack_0, ack => access_T_CP_0_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_202_Update/ack
      -- 
    ack_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_197_delayed_7_0_200_inst_ack_1, ack => access_T_CP_0_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	232 
    -- CP-element group 237: 	236 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (5) 
      -- CP-element group 237: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/word_access_start/$entry
      -- CP-element group 237: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/word_access_start/word_0/$entry
      -- CP-element group 237: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/word_access_start/word_0/rr
      -- 
    rr_873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(237), ack => ptr_deref_206_load_0_req_0); -- 
    access_T_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(232) & access_T_CP_0_elements(236) & access_T_CP_0_elements(239);
      gj_access_T_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	27 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (5) 
      -- CP-element group 238: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_update_start_
      -- CP-element group 238: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/word_access_complete/$entry
      -- CP-element group 238: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/word_access_complete/word_0/$entry
      -- CP-element group 238: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/word_access_complete/word_0/cr
      -- 
    cr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(238), ack => ptr_deref_206_load_0_req_1); -- 
    access_T_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(240);
      gj_access_T_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	227 
    -- CP-element group 239: 	234 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (5) 
      -- CP-element group 239: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/word_access_start/$exit
      -- CP-element group 239: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/word_access_start/word_0/$exit
      -- CP-element group 239: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Sample/word_access_start/word_0/ra
      -- 
    ra_874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_206_load_0_ack_0, ack => access_T_CP_0_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	313 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	110 
    -- CP-element group 240: 	238 
    -- CP-element group 240:  members (9) 
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/word_access_complete/$exit
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/word_access_complete/word_0/$exit
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/word_access_complete/word_0/ca
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/ptr_deref_206_Merge/$entry
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/ptr_deref_206_Merge/$exit
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/ptr_deref_206_Merge/merge_req
      -- CP-element group 240: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_206_Update/ptr_deref_206_Merge/merge_ack
      -- 
    ca_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_206_load_0_ack_1, ack => access_T_CP_0_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	35 
    -- CP-element group 241: 	225 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Sample/req
      -- 
    req_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(241), ack => W_fn1_203_delayed_13_0_208_inst_req_0); -- 
    access_T_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(35) & access_T_CP_0_elements(225) & access_T_CP_0_elements(243);
      gj_access_T_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	27 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_update_start_
      -- CP-element group 242: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Update/req
      -- 
    req_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(242), ack => W_fn1_203_delayed_13_0_208_inst_req_1); -- 
    access_T_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(244);
      gj_access_T_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	31 
    -- CP-element group 243: 	223 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Sample/ack
      -- 
    ack_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_203_delayed_13_0_208_inst_ack_0, ack => access_T_CP_0_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	313 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	110 
    -- CP-element group 244: 	242 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_210_Update/ack
      -- 
    ack_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_203_delayed_13_0_208_inst_ack_1, ack => access_T_CP_0_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	115 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Sample/req
      -- 
    req_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(245), ack => W_fetch_val1_205_delayed_13_0_211_inst_req_0); -- 
    access_T_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(115) & access_T_CP_0_elements(247);
      gj_access_T_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	27 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_update_start_
      -- CP-element group 246: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Update/req
      -- 
    req_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(246), ack => W_fetch_val1_205_delayed_13_0_211_inst_req_1); -- 
    access_T_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(248);
      gj_access_T_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	111 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Sample/ack
      -- 
    ack_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_205_delayed_13_0_211_inst_ack_0, ack => access_T_CP_0_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	313 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	110 
    -- CP-element group 248: 	246 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_213_Update/ack
      -- 
    ack_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_205_delayed_13_0_211_inst_ack_1, ack => access_T_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	115 
    -- CP-element group 249: 	35 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Sample/req
      -- 
    req_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(249), ack => WPIPE_input_pipe1_220_inst_req_0); -- 
    access_T_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(115) & access_T_CP_0_elements(35) & access_T_CP_0_elements(251);
      gj_access_T_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	111 
    -- CP-element group 250: 	31 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_update_start_
      -- CP-element group 250: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Sample/ack
      -- CP-element group 250: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Update/req
      -- 
    ack_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_220_inst_ack_0, ack => access_T_CP_0_elements(250)); -- 
    req_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(250), ack => WPIPE_input_pipe1_220_inst_req_1); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	313 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe1_220_Update/ack
      -- 
    ack_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_220_inst_ack_1, ack => access_T_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	96 
    -- CP-element group 252: 	170 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Sample/req
      -- 
    req_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(252), ack => W_continue_247_delayed_1_0_251_inst_req_0); -- 
    access_T_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(96) & access_T_CP_0_elements(170) & access_T_CP_0_elements(254);
      gj_access_T_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	265 
    -- CP-element group 253: 	273 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Update/req
      -- CP-element group 253: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_update_start_
      -- CP-element group 253: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Update/$entry
      -- 
    req_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(253), ack => W_continue_247_delayed_1_0_251_inst_req_1); -- 
    access_T_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(255) & access_T_CP_0_elements(265) & access_T_CP_0_elements(273);
      gj_access_T_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	92 
    -- CP-element group 254: 	166 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Sample/ack
      -- 
    ack_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_247_delayed_1_0_251_inst_ack_0, ack => access_T_CP_0_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	263 
    -- CP-element group 255: 	271 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Update/ack
      -- CP-element group 255: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_253_Update/$exit
      -- 
    ack_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_247_delayed_1_0_251_inst_ack_1, ack => access_T_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	260 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	261 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	261 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_request/req
      -- CP-element group 256: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_request/$entry
      -- 
    req_986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(256), ack => addr_of_272_final_reg_req_0); -- 
    access_T_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(260) & access_T_CP_0_elements(261);
      gj_access_T_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	24 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	262 
    -- CP-element group 257: 	269 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	262 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_complete/$entry
      -- CP-element group 257: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_complete/req
      -- CP-element group 257: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_update_start_
      -- 
    req_991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(257), ack => addr_of_272_final_reg_req_1); -- 
    access_T_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(262) & access_T_CP_0_elements(269);
      gj_access_T_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	24 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	261 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Update/req
      -- CP-element group 258: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_update_start
      -- 
    req_976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(258), ack => array_obj_ref_271_index_offset_req_1); -- 
    access_T_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(260) & access_T_CP_0_elements(261);
      gj_access_T_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	54 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	313 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	50 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_sample_complete
      -- 
    ack_972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_271_index_offset_ack_0, ack => access_T_CP_0_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	256 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260:  members (8) 
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_base_plus_offset/sum_rename_req
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_offset_calculated
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_base_plus_offset/sum_rename_ack
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_root_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_base_plus_offset/$exit
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_base_plus_offset/$entry
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_271_final_index_sum_regn_Update/$exit
      -- 
    ack_977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_271_index_offset_ack_1, ack => access_T_CP_0_elements(260)); -- 
    -- CP-element group 261:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	256 
    -- CP-element group 261: successors 
    -- CP-element group 261: marked-successors 
    -- CP-element group 261: 	256 
    -- CP-element group 261: 	258 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_request/ack
      -- CP-element group 261: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_request/$exit
      -- CP-element group 261: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_sample_completed_
      -- 
    ack_987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_272_final_reg_ack_0, ack => access_T_CP_0_elements(261)); -- 
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	267 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	257 
    -- CP-element group 262:  members (19) 
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_word_addrgen/$entry
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_word_addrgen/root_register_ack
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_complete/ack
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_word_addrgen/root_register_req
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_word_addrgen/$exit
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_plus_offset/sum_rename_ack
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_272_complete/$exit
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_plus_offset/sum_rename_req
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_plus_offset/$exit
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_plus_offset/$entry
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_addr_resize/base_resize_ack
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_addr_resize/base_resize_req
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_addr_resize/$exit
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_addr_resize/$entry
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_address_resized
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_root_address_calculated
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_word_address_calculated
      -- CP-element group 262: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_base_address_calculated
      -- 
    ack_992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_272_final_reg_ack_1, ack => access_T_CP_0_elements(262)); -- 
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	54 
    -- CP-element group 263: 	255 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Sample/req
      -- CP-element group 263: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_sample_start_
      -- 
    req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(263), ack => W_fn2_259_delayed_7_0_274_inst_req_0); -- 
    access_T_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(54) & access_T_CP_0_elements(255) & access_T_CP_0_elements(265);
      gj_access_T_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: 	269 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Update/req
      -- CP-element group 264: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_update_start_
      -- 
    req_1005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(264), ack => W_fn2_259_delayed_7_0_274_inst_req_1); -- 
    access_T_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(266) & access_T_CP_0_elements(269);
      gj_access_T_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: marked-successors 
    -- CP-element group 265: 	50 
    -- CP-element group 265: 	253 
    -- CP-element group 265: 	263 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_sample_completed_
      -- 
    ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_259_delayed_7_0_274_inst_ack_0, ack => access_T_CP_0_elements(265)); -- 
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_276_update_completed_
      -- 
    ack_1006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_259_delayed_7_0_274_inst_ack_1, ack => access_T_CP_0_elements(266)); -- 
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	266 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	269 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (5) 
      -- CP-element group 267: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/word_access_start/$entry
      -- CP-element group 267: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/word_access_start/word_0/rr
      -- CP-element group 267: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/word_access_start/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_sample_start_
      -- 
    rr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(267), ack => ptr_deref_280_load_0_req_0); -- 
    access_T_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(262) & access_T_CP_0_elements(266) & access_T_CP_0_elements(269);
      gj_access_T_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	27 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (5) 
      -- CP-element group 268: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/word_access_complete/$entry
      -- CP-element group 268: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/word_access_complete/word_0/cr
      -- CP-element group 268: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_update_start_
      -- CP-element group 268: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/word_access_complete/word_0/$entry
      -- 
    cr_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(268), ack => ptr_deref_280_load_0_req_1); -- 
    access_T_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(270);
      gj_access_T_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: marked-successors 
    -- CP-element group 269: 	257 
    -- CP-element group 269: 	264 
    -- CP-element group 269: 	267 
    -- CP-element group 269:  members (5) 
      -- CP-element group 269: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/word_access_start/word_0/ra
      -- CP-element group 269: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/word_access_start/word_0/$exit
      -- CP-element group 269: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/word_access_start/$exit
      -- CP-element group 269: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_sample_completed_
      -- 
    ra_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_280_load_0_ack_0, ack => access_T_CP_0_elements(269)); -- 
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	313 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	129 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (9) 
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/ptr_deref_280_Merge/merge_ack
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/word_access_complete/$exit
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/ptr_deref_280_Merge/merge_req
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/ptr_deref_280_Merge/$exit
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/ptr_deref_280_Merge/$entry
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/word_access_complete/word_0/ca
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_Update/word_access_complete/word_0/$exit
      -- CP-element group 270: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_280_update_completed_
      -- 
    ca_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_280_load_0_ack_1, ack => access_T_CP_0_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	54 
    -- CP-element group 271: 	255 
    -- CP-element group 271: marked-predecessors 
    -- CP-element group 271: 	273 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Sample/req
      -- CP-element group 271: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_sample_start_
      -- 
    req_1064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(271), ack => W_fn2_265_delayed_13_0_282_inst_req_0); -- 
    access_T_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(54) & access_T_CP_0_elements(255) & access_T_CP_0_elements(273);
      gj_access_T_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	27 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_update_start_
      -- CP-element group 272: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Update/req
      -- CP-element group 272: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Update/$entry
      -- 
    req_1069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(272), ack => W_fn2_265_delayed_13_0_282_inst_req_1); -- 
    access_T_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(274);
      gj_access_T_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273: marked-successors 
    -- CP-element group 273: 	50 
    -- CP-element group 273: 	253 
    -- CP-element group 273: 	271 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Sample/ack
      -- 
    ack_1065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_265_delayed_13_0_282_inst_ack_0, ack => access_T_CP_0_elements(273)); -- 
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	313 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	129 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_284_Update/$exit
      -- 
    ack_1070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_265_delayed_13_0_282_inst_ack_1, ack => access_T_CP_0_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	132 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	277 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Sample/req
      -- CP-element group 275: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Sample/$entry
      -- 
    req_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(275), ack => W_fetch_val2_267_delayed_13_0_285_inst_req_0); -- 
    access_T_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(132) & access_T_CP_0_elements(277);
      gj_access_T_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	27 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Update/req
      -- CP-element group 276: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Update/$entry
      -- CP-element group 276: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_update_start_
      -- 
    req_1083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(276), ack => W_fetch_val2_267_delayed_13_0_285_inst_req_1); -- 
    access_T_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(278);
      gj_access_T_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	130 
    -- CP-element group 277: 	275 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_sample_completed_
      -- 
    ack_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_267_delayed_13_0_285_inst_ack_0, ack => access_T_CP_0_elements(277)); -- 
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	313 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	129 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_287_update_completed_
      -- 
    ack_1084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_267_delayed_13_0_285_inst_ack_1, ack => access_T_CP_0_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	132 
    -- CP-element group 279: 	54 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Sample/req
      -- CP-element group 279: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_sample_start_
      -- 
    req_1092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(279), ack => WPIPE_input_pipe2_294_inst_req_0); -- 
    access_T_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(132) & access_T_CP_0_elements(54) & access_T_CP_0_elements(281);
      gj_access_T_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	130 
    -- CP-element group 280: 	50 
    -- CP-element group 280:  members (6) 
      -- CP-element group 280: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Update/req
      -- CP-element group 280: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Sample/ack
      -- CP-element group 280: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_update_start_
      -- CP-element group 280: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_sample_completed_
      -- 
    ack_1093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_294_inst_ack_0, ack => access_T_CP_0_elements(280)); -- 
    req_1097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(280), ack => WPIPE_input_pipe2_294_inst_req_1); -- 
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	313 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	279 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Update/ack
      -- CP-element group 281: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe2_294_update_completed_
      -- 
    ack_1098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_294_inst_ack_1, ack => access_T_CP_0_elements(281)); -- 
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	96 
    -- CP-element group 282: 	170 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	284 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Sample/req
      -- CP-element group 282: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_sample_start_
      -- 
    req_1106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(282), ack => W_continue_309_delayed_1_0_325_inst_req_0); -- 
    access_T_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(96) & access_T_CP_0_elements(170) & access_T_CP_0_elements(284);
      gj_access_T_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	285 
    -- CP-element group 283: 	295 
    -- CP-element group 283: 	303 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Update/req
      -- CP-element group 283: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_update_start_
      -- 
    req_1111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(283), ack => W_continue_309_delayed_1_0_325_inst_req_1); -- 
    access_T_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(285) & access_T_CP_0_elements(295) & access_T_CP_0_elements(303);
      gj_access_T_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	92 
    -- CP-element group 284: 	166 
    -- CP-element group 284: 	282 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_sample_completed_
      -- 
    ack_1107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_309_delayed_1_0_325_inst_ack_0, ack => access_T_CP_0_elements(284)); -- 
    -- CP-element group 285:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	293 
    -- CP-element group 285: 	301 
    -- CP-element group 285: marked-successors 
    -- CP-element group 285: 	283 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Update/ack
      -- CP-element group 285: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_327_update_completed_
      -- 
    ack_1112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_309_delayed_1_0_325_inst_ack_1, ack => access_T_CP_0_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	290 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	291 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	291 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_request/$entry
      -- CP-element group 286: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_request/req
      -- 
    req_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(286), ack => addr_of_351_final_reg_req_0); -- 
    access_T_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(290) & access_T_CP_0_elements(291);
      gj_access_T_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	24 
    -- CP-element group 287: marked-predecessors 
    -- CP-element group 287: 	292 
    -- CP-element group 287: 	299 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	292 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_complete/req
      -- CP-element group 287: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_complete/$entry
      -- CP-element group 287: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_update_start_
      -- 
    req_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(287), ack => addr_of_351_final_reg_req_1); -- 
    access_T_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(292) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	24 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	290 
    -- CP-element group 288: 	291 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_update_start
      -- CP-element group 288: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Update/req
      -- 
    req_1142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(288), ack => array_obj_ref_350_index_offset_req_1); -- 
    access_T_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(290) & access_T_CP_0_elements(291);
      gj_access_T_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	75 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	313 
    -- CP-element group 289: marked-successors 
    -- CP-element group 289: 	71 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_sample_complete
      -- 
    ack_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_350_index_offset_ack_0, ack => access_T_CP_0_elements(289)); -- 
    -- CP-element group 290:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	286 
    -- CP-element group 290: marked-successors 
    -- CP-element group 290: 	288 
    -- CP-element group 290:  members (8) 
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_base_plus_offset/sum_rename_ack
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_base_plus_offset/sum_rename_req
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_base_plus_offset/$exit
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_base_plus_offset/$entry
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_final_index_sum_regn_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_offset_calculated
      -- CP-element group 290: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/array_obj_ref_350_root_address_calculated
      -- 
    ack_1143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_350_index_offset_ack_1, ack => access_T_CP_0_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	286 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	286 
    -- CP-element group 291: 	288 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_request/ack
      -- CP-element group 291: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_request/$exit
      -- 
    ack_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_351_final_reg_ack_0, ack => access_T_CP_0_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	287 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	297 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	287 
    -- CP-element group 292:  members (19) 
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_addr_resize/base_resize_ack
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_addr_resize/base_resize_req
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_addr_resize/$exit
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_addr_resize/$entry
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_address_resized
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_root_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_complete/ack
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_word_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_word_addrgen/root_register_ack
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_plus_offset/sum_rename_ack
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_word_addrgen/root_register_req
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_word_addrgen/$exit
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_complete/$exit
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_plus_offset/sum_rename_req
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_plus_offset/$exit
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_base_plus_offset/$entry
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_word_addrgen/$entry
      -- CP-element group 292: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/addr_of_351_update_completed_
      -- 
    ack_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_351_final_reg_ack_1, ack => access_T_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	75 
    -- CP-element group 293: 	285 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_sample_start_
      -- 
    req_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(293), ack => W_fn3_326_delayed_7_0_353_inst_req_0); -- 
    access_T_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(285) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: 	299 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Update/req
      -- CP-element group 294: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_update_start_
      -- 
    req_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(294), ack => W_fn3_326_delayed_7_0_353_inst_req_1); -- 
    access_T_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(296) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	71 
    -- CP-element group 295: 	283 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_sample_completed_
      -- 
    ack_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_326_delayed_7_0_353_inst_ack_0, ack => access_T_CP_0_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_355_update_completed_
      -- 
    ack_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_326_delayed_7_0_353_inst_ack_1, ack => access_T_CP_0_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	292 
    -- CP-element group 297: 	296 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (5) 
      -- CP-element group 297: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/word_access_start/word_0/$entry
      -- CP-element group 297: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/word_access_start/$entry
      -- CP-element group 297: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/word_access_start/word_0/rr
      -- CP-element group 297: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_sample_start_
      -- 
    rr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(297), ack => ptr_deref_359_load_0_req_0); -- 
    access_T_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(292) & access_T_CP_0_elements(296) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	27 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (5) 
      -- CP-element group 298: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/word_access_complete/$entry
      -- CP-element group 298: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/word_access_complete/word_0/cr
      -- CP-element group 298: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/word_access_complete/word_0/$entry
      -- CP-element group 298: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_update_start_
      -- 
    cr_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(298), ack => ptr_deref_359_load_0_req_1); -- 
    access_T_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(300);
      gj_access_T_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	287 
    -- CP-element group 299: 	294 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (5) 
      -- CP-element group 299: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/word_access_start/$exit
      -- CP-element group 299: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/word_access_start/word_0/ra
      -- CP-element group 299: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Sample/word_access_start/word_0/$exit
      -- 
    ra_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_359_load_0_ack_0, ack => access_T_CP_0_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	313 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	146 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (9) 
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/ptr_deref_359_Merge/merge_ack
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/word_access_complete/word_0/ca
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/word_access_complete/word_0/$exit
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/word_access_complete/$exit
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/ptr_deref_359_Merge/merge_req
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/ptr_deref_359_Merge/$exit
      -- CP-element group 300: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/ptr_deref_359_Update/ptr_deref_359_Merge/$entry
      -- 
    ca_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_359_load_0_ack_1, ack => access_T_CP_0_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	75 
    -- CP-element group 301: 	285 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Sample/req
      -- CP-element group 301: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Sample/$entry
      -- 
    req_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(301), ack => W_fn3_332_delayed_13_0_361_inst_req_0); -- 
    access_T_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(285) & access_T_CP_0_elements(303);
      gj_access_T_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	27 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_update_start_
      -- CP-element group 302: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Update/req
      -- CP-element group 302: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Update/$entry
      -- 
    req_1235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(302), ack => W_fn3_332_delayed_13_0_361_inst_req_1); -- 
    access_T_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(304);
      gj_access_T_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	71 
    -- CP-element group 303: 	283 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Sample/ack
      -- 
    ack_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_332_delayed_13_0_361_inst_ack_0, ack => access_T_CP_0_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	313 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	146 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_363_Update/$exit
      -- 
    ack_1236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_332_delayed_13_0_361_inst_ack_1, ack => access_T_CP_0_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	151 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Sample/req
      -- 
    req_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(305), ack => W_fetch_val3_334_delayed_13_0_364_inst_req_0); -- 
    access_T_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(151) & access_T_CP_0_elements(307);
      gj_access_T_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	27 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_update_start_
      -- CP-element group 306: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Update/req
      -- 
    req_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(306), ack => W_fetch_val3_334_delayed_13_0_364_inst_req_1); -- 
    access_T_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	147 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Sample/ack
      -- 
    ack_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_334_delayed_13_0_364_inst_ack_0, ack => access_T_CP_0_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	313 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	146 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/assign_stmt_366_Update/ack
      -- 
    ack_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_334_delayed_13_0_364_inst_ack_1, ack => access_T_CP_0_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	75 
    -- CP-element group 309: 	151 
    -- CP-element group 309: 	170 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Sample/req
      -- 
    req_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(309), ack => WPIPE_input_pipe3_374_inst_req_0); -- 
    access_T_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(151) & access_T_CP_0_elements(170) & access_T_CP_0_elements(311);
      gj_access_T_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310: marked-successors 
    -- CP-element group 310: 	71 
    -- CP-element group 310: 	147 
    -- CP-element group 310: 	166 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_update_start_
      -- CP-element group 310: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Sample/ack
      -- CP-element group 310: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Update/req
      -- 
    ack_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_374_inst_ack_0, ack => access_T_CP_0_elements(310)); -- 
    req_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(310), ack => WPIPE_input_pipe3_374_inst_req_1); -- 
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	309 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/WPIPE_input_pipe3_374_Update/ack
      -- 
    ack_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_374_inst_ack_1, ack => access_T_CP_0_elements(311)); -- 
    -- CP-element group 312:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	24 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	25 
    -- CP-element group 312:  members (1) 
      -- CP-element group 312: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(312) is a control-delay.
    cp_element_312_delay: control_delay_element  generic map(name => " 312_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(24), ack => access_T_CP_0_elements(312), clk => clk, reset =>reset);
    -- CP-element group 313:  join  transition  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	27 
    -- CP-element group 313: 	229 
    -- CP-element group 313: 	240 
    -- CP-element group 313: 	244 
    -- CP-element group 313: 	248 
    -- CP-element group 313: 	251 
    -- CP-element group 313: 	259 
    -- CP-element group 313: 	270 
    -- CP-element group 313: 	274 
    -- CP-element group 313: 	278 
    -- CP-element group 313: 	281 
    -- CP-element group 313: 	289 
    -- CP-element group 313: 	300 
    -- CP-element group 313: 	304 
    -- CP-element group 313: 	308 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	21 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_28/do_while_stmt_81/do_while_stmt_81_loop_body/$exit
      -- 
    access_T_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(229) & access_T_CP_0_elements(240) & access_T_CP_0_elements(244) & access_T_CP_0_elements(248) & access_T_CP_0_elements(251) & access_T_CP_0_elements(259) & access_T_CP_0_elements(270) & access_T_CP_0_elements(274) & access_T_CP_0_elements(278) & access_T_CP_0_elements(281) & access_T_CP_0_elements(289) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304) & access_T_CP_0_elements(308) & access_T_CP_0_elements(311);
      gj_access_T_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	20 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (2) 
      -- CP-element group 314: 	 branch_block_stmt_28/do_while_stmt_81/loop_exit/$exit
      -- CP-element group 314: 	 branch_block_stmt_28/do_while_stmt_81/loop_exit/ack
      -- 
    ack_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_81_branch_ack_0, ack => access_T_CP_0_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	20 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_28/do_while_stmt_81/loop_taken/$exit
      -- CP-element group 315: 	 branch_block_stmt_28/do_while_stmt_81/loop_taken/ack
      -- 
    ack_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_81_branch_ack_1, ack => access_T_CP_0_elements(315)); -- 
    -- CP-element group 316:  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	18 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	1 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_28/do_while_stmt_81/$exit
      -- 
    access_T_CP_0_elements(316) <= access_T_CP_0_elements(18);
    access_T_do_while_stmt_81_terminator_1274: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_81_terminator_1274", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(21),loop_continue => access_T_CP_0_elements(315),loop_terminate => access_T_CP_0_elements(314),loop_back => access_T_CP_0_elements(19),loop_exit => access_T_CP_0_elements(18),clk => clk, reset => reset); -- 
    phi_stmt_83_phi_seq_320_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(38);
      access_T_CP_0_elements(41)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(41);
      access_T_CP_0_elements(42)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(43);
      access_T_CP_0_elements(39) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(36);
      access_T_CP_0_elements(45)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(46)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(48);
      access_T_CP_0_elements(37) <= phi_mux_reqs(1);
      phi_stmt_83_phi_seq_320 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_83_phi_seq_320") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(32), 
          phi_sample_ack => access_T_CP_0_elements(33), 
          phi_update_req => access_T_CP_0_elements(34), 
          phi_update_ack => access_T_CP_0_elements(35), 
          phi_mux_ack => access_T_CP_0_elements(40), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_88_phi_seq_374_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(57);
      access_T_CP_0_elements(60)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(64);
      access_T_CP_0_elements(61)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(65);
      access_T_CP_0_elements(58) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(55);
      access_T_CP_0_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(68);
      access_T_CP_0_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(69);
      access_T_CP_0_elements(56) <= phi_mux_reqs(1);
      phi_stmt_88_phi_seq_374 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_88_phi_seq_374") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(51), 
          phi_sample_ack => access_T_CP_0_elements(52), 
          phi_update_req => access_T_CP_0_elements(53), 
          phi_update_ack => access_T_CP_0_elements(54), 
          phi_mux_ack => access_T_CP_0_elements(59), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_93_phi_seq_428_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(85);
      access_T_CP_0_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(86);
      access_T_CP_0_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(76);
      access_T_CP_0_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(77) <= phi_mux_reqs(1);
      phi_stmt_93_phi_seq_428 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_93_phi_seq_428") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(72), 
          phi_sample_ack => access_T_CP_0_elements(73), 
          phi_update_req => access_T_CP_0_elements(74), 
          phi_update_ack => access_T_CP_0_elements(75), 
          phi_mux_ack => access_T_CP_0_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_98_phi_seq_472_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(102)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(102);
      access_T_CP_0_elements(103)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(100) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(97);
      access_T_CP_0_elements(106)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(108);
      access_T_CP_0_elements(107)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(109);
      access_T_CP_0_elements(98) <= phi_mux_reqs(1);
      phi_stmt_98_phi_seq_472 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_98_phi_seq_472") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(93), 
          phi_sample_ack => access_T_CP_0_elements(94), 
          phi_update_req => access_T_CP_0_elements(95), 
          phi_update_ack => access_T_CP_0_elements(96), 
          phi_mux_ack => access_T_CP_0_elements(101), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_103_phi_seq_526_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(121)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(123);
      access_T_CP_0_elements(122)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(124);
      access_T_CP_0_elements(119) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(125)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(126)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(128);
      access_T_CP_0_elements(117) <= phi_mux_reqs(1);
      phi_stmt_103_phi_seq_526 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_103_phi_seq_526") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(112), 
          phi_sample_ack => access_T_CP_0_elements(113), 
          phi_update_req => access_T_CP_0_elements(114), 
          phi_update_ack => access_T_CP_0_elements(115), 
          phi_mux_ack => access_T_CP_0_elements(120), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_107_phi_seq_580_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(138)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(140);
      access_T_CP_0_elements(139)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(141);
      access_T_CP_0_elements(136) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(133);
      access_T_CP_0_elements(142)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(144);
      access_T_CP_0_elements(143)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(145);
      access_T_CP_0_elements(134) <= phi_mux_reqs(1);
      phi_stmt_107_phi_seq_580 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_107_phi_seq_580") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(26), 
          phi_sample_ack => access_T_CP_0_elements(131), 
          phi_update_req => access_T_CP_0_elements(28), 
          phi_update_ack => access_T_CP_0_elements(132), 
          phi_mux_ack => access_T_CP_0_elements(137), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_111_phi_seq_634_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(154);
      access_T_CP_0_elements(157)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(159);
      access_T_CP_0_elements(158)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(160);
      access_T_CP_0_elements(155) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(152);
      access_T_CP_0_elements(161)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(163);
      access_T_CP_0_elements(162)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(164);
      access_T_CP_0_elements(153) <= phi_mux_reqs(1);
      phi_stmt_111_phi_seq_634 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_111_phi_seq_634") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(148), 
          phi_sample_ack => access_T_CP_0_elements(149), 
          phi_update_req => access_T_CP_0_elements(150), 
          phi_update_ack => access_T_CP_0_elements(151), 
          phi_mux_ack => access_T_CP_0_elements(156), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_115_phi_seq_678_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(173);
      access_T_CP_0_elements(176)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(176);
      access_T_CP_0_elements(177)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(178);
      access_T_CP_0_elements(174) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(171);
      access_T_CP_0_elements(180)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(182);
      access_T_CP_0_elements(181)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(183);
      access_T_CP_0_elements(172) <= phi_mux_reqs(1);
      phi_stmt_115_phi_seq_678 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_115_phi_seq_678") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(167), 
          phi_sample_ack => access_T_CP_0_elements(168), 
          phi_update_req => access_T_CP_0_elements(169), 
          phi_update_ack => access_T_CP_0_elements(170), 
          phi_mux_ack => access_T_CP_0_elements(175), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_120_phi_seq_722_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(192);
      access_T_CP_0_elements(195)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(195);
      access_T_CP_0_elements(196)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(197);
      access_T_CP_0_elements(193) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(190);
      access_T_CP_0_elements(199)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(201);
      access_T_CP_0_elements(200)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(202);
      access_T_CP_0_elements(191) <= phi_mux_reqs(1);
      phi_stmt_120_phi_seq_722 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_120_phi_seq_722") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(186), 
          phi_sample_ack => access_T_CP_0_elements(187), 
          phi_update_req => access_T_CP_0_elements(188), 
          phi_update_ack => access_T_CP_0_elements(189), 
          phi_mux_ack => access_T_CP_0_elements(194), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_125_phi_seq_766_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(211);
      access_T_CP_0_elements(214)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(214);
      access_T_CP_0_elements(215)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(216);
      access_T_CP_0_elements(212) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(209);
      access_T_CP_0_elements(218)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(220);
      access_T_CP_0_elements(219)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(221);
      access_T_CP_0_elements(210) <= phi_mux_reqs(1);
      phi_stmt_125_phi_seq_766 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_125_phi_seq_766") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(205), 
          phi_sample_ack => access_T_CP_0_elements(206), 
          phi_update_req => access_T_CP_0_elements(207), 
          phi_update_ack => access_T_CP_0_elements(208), 
          phi_mux_ack => access_T_CP_0_elements(213), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_272_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(22);
        preds(1)  <= access_T_CP_0_elements(23);
        entry_tmerge_272 : transition_merge -- 
          generic map(name => " entry_tmerge_272")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(24));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_168_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_316_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_141_wire : std_logic_vector(31 downto 0);
    signal AND_u64_u64_153_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_227_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_301_wire : std_logic_vector(63 downto 0);
    signal LSHR_u32_u32_58_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_72_wire : std_logic_vector(31 downto 0);
    signal LSHR_u64_u64_161_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_183_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_186_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_196_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_196_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_196_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_235_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_257_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_260_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_270_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_270_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_270_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_309_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_331_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_334_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_349_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_349_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_349_wire : std_logic_vector(63 downto 0);
    signal MUL_u16_u16_33_wire : std_logic_vector(15 downto 0);
    signal NEQ_u64_u1_187_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_261_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_335_wire : std_logic_vector(0 downto 0);
    signal SUB_u64_u64_154_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_228_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_302_wire : std_logic_vector(63 downto 0);
    signal address1_83 : std_logic_vector(63 downto 0);
    signal address2_88 : std_logic_vector(63 downto 0);
    signal address3_93 : std_logic_vector(63 downto 0);
    signal array_obj_ref_197_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_197_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_197_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_197_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_197_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_197_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_271_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_271_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_271_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_271_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_271_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_271_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_74_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_74_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_74_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_74_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_74_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_74_root_address : std_logic_vector(13 downto 0);
    signal continue_148 : std_logic_vector(0 downto 0);
    signal continue_185_delayed_1_0_179 : std_logic_vector(0 downto 0);
    signal continue_247_delayed_1_0_253 : std_logic_vector(0 downto 0);
    signal continue_309_delayed_1_0_327 : std_logic_vector(0 downto 0);
    signal fetch_add1_48 : std_logic_vector(31 downto 0);
    signal fetch_add2_62 : std_logic_vector(31 downto 0);
    signal fetch_add3_76 : std_logic_vector(31 downto 0);
    signal fetch_addr1_199 : std_logic_vector(31 downto 0);
    signal fetch_addr2_273 : std_logic_vector(31 downto 0);
    signal fetch_addr3_352 : std_logic_vector(31 downto 0);
    signal fetch_val1_103 : std_logic_vector(63 downto 0);
    signal fetch_val1_205_delayed_13_0_213 : std_logic_vector(63 downto 0);
    signal fetch_val2_107 : std_logic_vector(63 downto 0);
    signal fetch_val2_267_delayed_13_0_287 : std_logic_vector(63 downto 0);
    signal fetch_val3_111 : std_logic_vector(63 downto 0);
    signal fetch_val3_334_delayed_13_0_366 : std_logic_vector(63 downto 0);
    signal fn1_190 : std_logic_vector(0 downto 0);
    signal fn1_197_delayed_7_0_202 : std_logic_vector(0 downto 0);
    signal fn1_203_delayed_13_0_210 : std_logic_vector(0 downto 0);
    signal fn2_259_delayed_7_0_276 : std_logic_vector(0 downto 0);
    signal fn2_264 : std_logic_vector(0 downto 0);
    signal fn2_265_delayed_13_0_284 : std_logic_vector(0 downto 0);
    signal fn3_326_delayed_7_0_355 : std_logic_vector(0 downto 0);
    signal fn3_332_delayed_13_0_363 : std_logic_vector(0 downto 0);
    signal fn3_338 : std_logic_vector(0 downto 0);
    signal fv1_207 : std_logic_vector(63 downto 0);
    signal fv2_281 : std_logic_vector(63 downto 0);
    signal fv3_360 : std_logic_vector(63 downto 0);
    signal konst_138_wire_constant : std_logic_vector(31 downto 0);
    signal konst_140_wire_constant : std_logic_vector(31 downto 0);
    signal konst_150_wire_constant : std_logic_vector(63 downto 0);
    signal konst_152_wire_constant : std_logic_vector(63 downto 0);
    signal konst_155_wire_constant : std_logic_vector(63 downto 0);
    signal konst_167_wire_constant : std_logic_vector(15 downto 0);
    signal konst_174_wire_constant : std_logic_vector(63 downto 0);
    signal konst_182_wire_constant : std_logic_vector(63 downto 0);
    signal konst_185_wire_constant : std_logic_vector(63 downto 0);
    signal konst_195_wire_constant : std_logic_vector(63 downto 0);
    signal konst_224_wire_constant : std_logic_vector(63 downto 0);
    signal konst_226_wire_constant : std_logic_vector(63 downto 0);
    signal konst_229_wire_constant : std_logic_vector(63 downto 0);
    signal konst_241_wire_constant : std_logic_vector(15 downto 0);
    signal konst_248_wire_constant : std_logic_vector(63 downto 0);
    signal konst_256_wire_constant : std_logic_vector(63 downto 0);
    signal konst_259_wire_constant : std_logic_vector(63 downto 0);
    signal konst_269_wire_constant : std_logic_vector(63 downto 0);
    signal konst_298_wire_constant : std_logic_vector(63 downto 0);
    signal konst_300_wire_constant : std_logic_vector(63 downto 0);
    signal konst_303_wire_constant : std_logic_vector(63 downto 0);
    signal konst_315_wire_constant : std_logic_vector(15 downto 0);
    signal konst_322_wire_constant : std_logic_vector(63 downto 0);
    signal konst_330_wire_constant : std_logic_vector(63 downto 0);
    signal konst_333_wire_constant : std_logic_vector(63 downto 0);
    signal konst_348_wire_constant : std_logic_vector(63 downto 0);
    signal konst_38_wire_constant : std_logic_vector(31 downto 0);
    signal konst_57_wire_constant : std_logic_vector(31 downto 0);
    signal konst_71_wire_constant : std_logic_vector(31 downto 0);
    signal m2_factor_40 : std_logic_vector(31 downto 0);
    signal m_factor_35 : std_logic_vector(31 downto 0);
    signal my_fetch1_52 : std_logic_vector(63 downto 0);
    signal my_fetch1_52_105_buffered : std_logic_vector(63 downto 0);
    signal my_fetch2_66 : std_logic_vector(63 downto 0);
    signal my_fetch2_66_109_buffered : std_logic_vector(63 downto 0);
    signal my_fetch3_80 : std_logic_vector(63 downto 0);
    signal my_fetch3_80_113_buffered : std_logic_vector(63 downto 0);
    signal my_num1_157 : std_logic_vector(63 downto 0);
    signal my_num2_231 : std_logic_vector(63 downto 0);
    signal my_num3_305 : std_logic_vector(63 downto 0);
    signal mycounter_98 : std_logic_vector(31 downto 0);
    signal n_address1_176 : std_logic_vector(63 downto 0);
    signal n_address1_176_87_buffered : std_logic_vector(63 downto 0);
    signal n_address2_250 : std_logic_vector(63 downto 0);
    signal n_address2_250_92_buffered : std_logic_vector(63 downto 0);
    signal n_address3_324 : std_logic_vector(63 downto 0);
    signal n_address3_324_97_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val1_219 : std_logic_vector(63 downto 0);
    signal n_fetch_val1_219_106_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val2_293 : std_logic_vector(63 downto 0);
    signal n_fetch_val2_293_110_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val3_372 : std_logic_vector(63 downto 0);
    signal n_fetch_val3_372_114_buffered : std_logic_vector(63 downto 0);
    signal n_mycounter_143 : std_logic_vector(31 downto 0);
    signal n_mycounter_143_102_buffered : std_logic_vector(31 downto 0);
    signal n_row1_171 : std_logic_vector(15 downto 0);
    signal n_row1_171_119_buffered : std_logic_vector(15 downto 0);
    signal n_row2_245 : std_logic_vector(15 downto 0);
    signal n_row2_245_124_buffered : std_logic_vector(15 downto 0);
    signal n_row3_319 : std_logic_vector(15 downto 0);
    signal n_row3_319_129_buffered : std_logic_vector(15 downto 0);
    signal next_row_135 : std_logic_vector(0 downto 0);
    signal ptr_deref_206_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_206_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_206_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_206_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_206_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_280_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_280_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_280_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_280_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_280_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_359_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_359_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_359_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_359_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_359_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_51_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_51_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_51_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_51_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_51_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_65_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_65_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_65_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_65_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_65_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_79_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_79_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_79_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_79_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_79_word_offset_0 : std_logic_vector(13 downto 0);
    signal row1_115 : std_logic_vector(15 downto 0);
    signal row2_120 : std_logic_vector(15 downto 0);
    signal row3_125 : std_logic_vector(15 downto 0);
    signal send_now3_343 : std_logic_vector(0 downto 0);
    signal type_cast_101_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_123_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_128_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_59_resized : std_logic_vector(13 downto 0);
    signal type_cast_59_scaled : std_logic_vector(13 downto 0);
    signal type_cast_59_wire : std_logic_vector(63 downto 0);
    signal type_cast_73_resized : std_logic_vector(13 downto 0);
    signal type_cast_73_scaled : std_logic_vector(13 downto 0);
    signal type_cast_73_wire : std_logic_vector(63 downto 0);
    signal type_cast_86_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_91_wire : std_logic_vector(63 downto 0);
    signal type_cast_96_wire : std_logic_vector(63 downto 0);
    signal var_val1_163 : std_logic_vector(15 downto 0);
    signal var_val2_237 : std_logic_vector(15 downto 0);
    signal var_val3_311 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_197_constant_part_of_offset <= "00000000000000";
    array_obj_ref_197_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_197_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_197_resized_base_address <= "00000000000000";
    array_obj_ref_271_constant_part_of_offset <= "00000000000000";
    array_obj_ref_271_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_271_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_271_resized_base_address <= "00000000000000";
    array_obj_ref_350_constant_part_of_offset <= "00000000000000";
    array_obj_ref_350_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_350_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_350_resized_base_address <= "00000000000000";
    array_obj_ref_60_constant_part_of_offset <= "00000000000000";
    array_obj_ref_60_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_60_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_60_resized_base_address <= "00000000000000";
    array_obj_ref_74_constant_part_of_offset <= "00000000000000";
    array_obj_ref_74_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_74_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_74_resized_base_address <= "00000000000000";
    fetch_add1_48 <= "00000000000000000000000000000000";
    konst_138_wire_constant <= "00000000000000000000000000000001";
    konst_140_wire_constant <= "00000000000000000000000000000001";
    konst_150_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_152_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_155_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_167_wire_constant <= "0000000000000001";
    konst_174_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_182_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_185_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_224_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_226_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_229_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_241_wire_constant <= "0000000000000001";
    konst_248_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_256_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_259_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_269_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_298_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_300_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_303_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_315_wire_constant <= "0000000000000001";
    konst_322_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_330_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_333_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_348_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_38_wire_constant <= "00000000000000000000000000000001";
    konst_57_wire_constant <= "00000000000000000000000000000010";
    konst_71_wire_constant <= "00000000000000000000000000000001";
    ptr_deref_206_word_offset_0 <= "00000000000000";
    ptr_deref_280_word_offset_0 <= "00000000000000";
    ptr_deref_359_word_offset_0 <= "00000000000000";
    ptr_deref_51_word_offset_0 <= "00000000000000";
    ptr_deref_65_word_offset_0 <= "00000000000000";
    ptr_deref_79_word_offset_0 <= "00000000000000";
    type_cast_101_wire_constant <= "00000000000000000000000000000001";
    type_cast_118_wire_constant <= "0000000000000000";
    type_cast_123_wire_constant <= "0000000000000001";
    type_cast_128_wire_constant <= "0000000000000010";
    type_cast_86_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_103: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch1_52_105_buffered & n_fetch_val1_219_106_buffered;
      req <= phi_stmt_103_req_0 & phi_stmt_103_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_103",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_103_ack_0,
          idata => idata,
          odata => fetch_val1_103,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_103
    phi_stmt_107: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch2_66_109_buffered & n_fetch_val2_293_110_buffered;
      req <= phi_stmt_107_req_0 & phi_stmt_107_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_107",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_107_ack_0,
          idata => idata,
          odata => fetch_val2_107,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_107
    phi_stmt_111: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch3_80_113_buffered & n_fetch_val3_372_114_buffered;
      req <= phi_stmt_111_req_0 & phi_stmt_111_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_111",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_111_ack_0,
          idata => idata,
          odata => fetch_val3_111,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_111
    phi_stmt_115: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_118_wire_constant & n_row1_171_119_buffered;
      req <= phi_stmt_115_req_0 & phi_stmt_115_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_115",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_115_ack_0,
          idata => idata,
          odata => row1_115,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_115
    phi_stmt_120: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_123_wire_constant & n_row2_245_124_buffered;
      req <= phi_stmt_120_req_0 & phi_stmt_120_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_120",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_120_ack_0,
          idata => idata,
          odata => row2_120,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_120
    phi_stmt_125: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_128_wire_constant & n_row3_319_129_buffered;
      req <= phi_stmt_125_req_0 & phi_stmt_125_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_125",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_125_ack_0,
          idata => idata,
          odata => row3_125,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_125
    phi_stmt_83: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_86_wire_constant & n_address1_176_87_buffered;
      req <= phi_stmt_83_req_0 & phi_stmt_83_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_83",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_83_ack_0,
          idata => idata,
          odata => address1_83,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_83
    phi_stmt_88: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_91_wire & n_address2_250_92_buffered;
      req <= phi_stmt_88_req_0 & phi_stmt_88_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_88",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_88_ack_0,
          idata => idata,
          odata => address2_88,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_88
    phi_stmt_93: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_96_wire & n_address3_324_97_buffered;
      req <= phi_stmt_93_req_0 & phi_stmt_93_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_93",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_93_ack_0,
          idata => idata,
          odata => address3_93,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_93
    phi_stmt_98: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_101_wire_constant & n_mycounter_143_102_buffered;
      req <= phi_stmt_98_req_0 & phi_stmt_98_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_98",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_98_ack_0,
          idata => idata,
          odata => mycounter_98,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_98
    -- flow-through select operator MUX_142_inst
    n_mycounter_143 <= konst_138_wire_constant when (next_row_135(0) /=  '0') else ADD_u32_u32_141_wire;
    -- flow-through select operator MUX_170_inst
    n_row1_171 <= ADD_u16_u16_168_wire when (next_row_135(0) /=  '0') else row1_115;
    -- flow-through select operator MUX_218_inst
    n_fetch_val1_219 <= fv1_207 when (fn1_203_delayed_13_0_210(0) /=  '0') else fetch_val1_205_delayed_13_0_213;
    -- flow-through select operator MUX_244_inst
    n_row2_245 <= ADD_u16_u16_242_wire when (next_row_135(0) /=  '0') else row2_120;
    -- flow-through select operator MUX_292_inst
    n_fetch_val2_293 <= fv2_281 when (fn2_265_delayed_13_0_284(0) /=  '0') else fetch_val2_267_delayed_13_0_287;
    -- flow-through select operator MUX_318_inst
    n_row3_319 <= ADD_u16_u16_316_wire when (next_row_135(0) /=  '0') else row3_125;
    -- flow-through select operator MUX_371_inst
    n_fetch_val3_372 <= fv3_360 when (fn3_332_delayed_13_0_363(0) /=  '0') else fetch_val3_334_delayed_13_0_366;
    W_continue_185_delayed_1_0_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_continue_185_delayed_1_0_177_inst_req_0;
      W_continue_185_delayed_1_0_177_inst_ack_0<= wack(0);
      rreq(0) <= W_continue_185_delayed_1_0_177_inst_req_1;
      W_continue_185_delayed_1_0_177_inst_ack_1<= rack(0);
      W_continue_185_delayed_1_0_177_inst : InterlockBuffer generic map ( -- 
        name => "W_continue_185_delayed_1_0_177_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => continue_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => continue_185_delayed_1_0_179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_continue_247_delayed_1_0_251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_continue_247_delayed_1_0_251_inst_req_0;
      W_continue_247_delayed_1_0_251_inst_ack_0<= wack(0);
      rreq(0) <= W_continue_247_delayed_1_0_251_inst_req_1;
      W_continue_247_delayed_1_0_251_inst_ack_1<= rack(0);
      W_continue_247_delayed_1_0_251_inst : InterlockBuffer generic map ( -- 
        name => "W_continue_247_delayed_1_0_251_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => continue_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => continue_247_delayed_1_0_253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_continue_309_delayed_1_0_325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_continue_309_delayed_1_0_325_inst_req_0;
      W_continue_309_delayed_1_0_325_inst_ack_0<= wack(0);
      rreq(0) <= W_continue_309_delayed_1_0_325_inst_req_1;
      W_continue_309_delayed_1_0_325_inst_ack_1<= rack(0);
      W_continue_309_delayed_1_0_325_inst : InterlockBuffer generic map ( -- 
        name => "W_continue_309_delayed_1_0_325_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => continue_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => continue_309_delayed_1_0_327,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val1_205_delayed_13_0_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val1_205_delayed_13_0_211_inst_req_0;
      W_fetch_val1_205_delayed_13_0_211_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val1_205_delayed_13_0_211_inst_req_1;
      W_fetch_val1_205_delayed_13_0_211_inst_ack_1<= rack(0);
      W_fetch_val1_205_delayed_13_0_211_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val1_205_delayed_13_0_211_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val1_103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val1_205_delayed_13_0_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val2_267_delayed_13_0_285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val2_267_delayed_13_0_285_inst_req_0;
      W_fetch_val2_267_delayed_13_0_285_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val2_267_delayed_13_0_285_inst_req_1;
      W_fetch_val2_267_delayed_13_0_285_inst_ack_1<= rack(0);
      W_fetch_val2_267_delayed_13_0_285_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val2_267_delayed_13_0_285_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val2_107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val2_267_delayed_13_0_287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val3_334_delayed_13_0_364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val3_334_delayed_13_0_364_inst_req_0;
      W_fetch_val3_334_delayed_13_0_364_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val3_334_delayed_13_0_364_inst_req_1;
      W_fetch_val3_334_delayed_13_0_364_inst_ack_1<= rack(0);
      W_fetch_val3_334_delayed_13_0_364_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val3_334_delayed_13_0_364_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val3_111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val3_334_delayed_13_0_366,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_197_delayed_7_0_200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_197_delayed_7_0_200_inst_req_0;
      W_fn1_197_delayed_7_0_200_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_197_delayed_7_0_200_inst_req_1;
      W_fn1_197_delayed_7_0_200_inst_ack_1<= rack(0);
      W_fn1_197_delayed_7_0_200_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_197_delayed_7_0_200_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_197_delayed_7_0_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_203_delayed_13_0_208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_203_delayed_13_0_208_inst_req_0;
      W_fn1_203_delayed_13_0_208_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_203_delayed_13_0_208_inst_req_1;
      W_fn1_203_delayed_13_0_208_inst_ack_1<= rack(0);
      W_fn1_203_delayed_13_0_208_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_203_delayed_13_0_208_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_203_delayed_13_0_210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_259_delayed_7_0_274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_259_delayed_7_0_274_inst_req_0;
      W_fn2_259_delayed_7_0_274_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_259_delayed_7_0_274_inst_req_1;
      W_fn2_259_delayed_7_0_274_inst_ack_1<= rack(0);
      W_fn2_259_delayed_7_0_274_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_259_delayed_7_0_274_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_259_delayed_7_0_276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_265_delayed_13_0_282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_265_delayed_13_0_282_inst_req_0;
      W_fn2_265_delayed_13_0_282_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_265_delayed_13_0_282_inst_req_1;
      W_fn2_265_delayed_13_0_282_inst_ack_1<= rack(0);
      W_fn2_265_delayed_13_0_282_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_265_delayed_13_0_282_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_265_delayed_13_0_284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_326_delayed_7_0_353_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_326_delayed_7_0_353_inst_req_0;
      W_fn3_326_delayed_7_0_353_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_326_delayed_7_0_353_inst_req_1;
      W_fn3_326_delayed_7_0_353_inst_ack_1<= rack(0);
      W_fn3_326_delayed_7_0_353_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_326_delayed_7_0_353_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_326_delayed_7_0_355,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_332_delayed_13_0_361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_332_delayed_13_0_361_inst_req_0;
      W_fn3_332_delayed_13_0_361_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_332_delayed_13_0_361_inst_req_1;
      W_fn3_332_delayed_13_0_361_inst_ack_1<= rack(0);
      W_fn3_332_delayed_13_0_361_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_332_delayed_13_0_361_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_332_delayed_13_0_363,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_198_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_198_final_reg_req_0;
      addr_of_198_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_198_final_reg_req_1;
      addr_of_198_final_reg_ack_1<= rack(0);
      addr_of_198_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_198_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_197_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_272_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_272_final_reg_req_0;
      addr_of_272_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_272_final_reg_req_1;
      addr_of_272_final_reg_ack_1<= rack(0);
      addr_of_272_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_272_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_271_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_273,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_351_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_351_final_reg_req_0;
      addr_of_351_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_351_final_reg_req_1;
      addr_of_351_final_reg_ack_1<= rack(0);
      addr_of_351_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_351_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_350_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr3_352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_61_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_61_final_reg_req_0;
      addr_of_61_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_61_final_reg_req_1;
      addr_of_61_final_reg_ack_1<= rack(0);
      addr_of_61_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_61_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_60_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add2_62,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_75_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_75_final_reg_req_0;
      addr_of_75_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_75_final_reg_req_1;
      addr_of_75_final_reg_ack_1<= rack(0);
      addr_of_75_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_75_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_74_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add3_76,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch1_52_105_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch1_52_105_buf_req_0;
      my_fetch1_52_105_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch1_52_105_buf_req_1;
      my_fetch1_52_105_buf_ack_1<= rack(0);
      my_fetch1_52_105_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch1_52_105_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch1_52,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch1_52_105_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch2_66_109_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch2_66_109_buf_req_0;
      my_fetch2_66_109_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch2_66_109_buf_req_1;
      my_fetch2_66_109_buf_ack_1<= rack(0);
      my_fetch2_66_109_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch2_66_109_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch2_66,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch2_66_109_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch3_80_113_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch3_80_113_buf_req_0;
      my_fetch3_80_113_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch3_80_113_buf_req_1;
      my_fetch3_80_113_buf_ack_1<= rack(0);
      my_fetch3_80_113_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch3_80_113_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch3_80,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch3_80_113_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_176_87_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_176_87_buf_req_0;
      n_address1_176_87_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_176_87_buf_req_1;
      n_address1_176_87_buf_ack_1<= rack(0);
      n_address1_176_87_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_176_87_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_176_87_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_250_92_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_250_92_buf_req_0;
      n_address2_250_92_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_250_92_buf_req_1;
      n_address2_250_92_buf_ack_1<= rack(0);
      n_address2_250_92_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_250_92_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_250_92_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address3_324_97_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address3_324_97_buf_req_0;
      n_address3_324_97_buf_ack_0<= wack(0);
      rreq(0) <= n_address3_324_97_buf_req_1;
      n_address3_324_97_buf_ack_1<= rack(0);
      n_address3_324_97_buf : InterlockBuffer generic map ( -- 
        name => "n_address3_324_97_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address3_324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address3_324_97_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val1_219_106_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val1_219_106_buf_req_0;
      n_fetch_val1_219_106_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val1_219_106_buf_req_1;
      n_fetch_val1_219_106_buf_ack_1<= rack(0);
      n_fetch_val1_219_106_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val1_219_106_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val1_219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val1_219_106_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val2_293_110_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val2_293_110_buf_req_0;
      n_fetch_val2_293_110_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val2_293_110_buf_req_1;
      n_fetch_val2_293_110_buf_ack_1<= rack(0);
      n_fetch_val2_293_110_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val2_293_110_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val2_293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val2_293_110_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val3_372_114_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val3_372_114_buf_req_0;
      n_fetch_val3_372_114_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val3_372_114_buf_req_1;
      n_fetch_val3_372_114_buf_ack_1<= rack(0);
      n_fetch_val3_372_114_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val3_372_114_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val3_372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val3_372_114_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter_143_102_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter_143_102_buf_req_0;
      n_mycounter_143_102_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter_143_102_buf_req_1;
      n_mycounter_143_102_buf_ack_1<= rack(0);
      n_mycounter_143_102_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter_143_102_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter_143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter_143_102_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row1_171_119_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row1_171_119_buf_req_0;
      n_row1_171_119_buf_ack_0<= wack(0);
      rreq(0) <= n_row1_171_119_buf_req_1;
      n_row1_171_119_buf_ack_1<= rack(0);
      n_row1_171_119_buf : InterlockBuffer generic map ( -- 
        name => "n_row1_171_119_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row1_171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row1_171_119_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row2_245_124_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row2_245_124_buf_req_0;
      n_row2_245_124_buf_ack_0<= wack(0);
      rreq(0) <= n_row2_245_124_buf_req_1;
      n_row2_245_124_buf_ack_1<= rack(0);
      n_row2_245_124_buf : InterlockBuffer generic map ( -- 
        name => "n_row2_245_124_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row2_245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row2_245_124_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row3_319_129_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row3_319_129_buf_req_0;
      n_row3_319_129_buf_ack_0<= wack(0);
      rreq(0) <= n_row3_319_129_buf_req_1;
      n_row3_319_129_buf_ack_1<= rack(0);
      n_row3_319_129_buf : InterlockBuffer generic map ( -- 
        name => "n_row3_319_129_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row3_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row3_319_129_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_162_inst
    process(LSHR_u64_u64_161_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_161_wire(15 downto 0);
      var_val1_163 <= tmp_var; -- 
    end process;
    -- interlock type_cast_236_inst
    process(LSHR_u64_u64_235_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_235_wire(15 downto 0);
      var_val2_237 <= tmp_var; -- 
    end process;
    -- interlock type_cast_310_inst
    process(LSHR_u64_u64_309_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_309_wire(15 downto 0);
      var_val3_311 <= tmp_var; -- 
    end process;
    -- interlock type_cast_34_inst
    process(MUL_u16_u16_33_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_33_wire(15 downto 0);
      m_factor_35 <= tmp_var; -- 
    end process;
    -- interlock type_cast_59_inst
    process(LSHR_u32_u32_58_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_58_wire(31 downto 0);
      type_cast_59_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_73_inst
    process(LSHR_u32_u32_72_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_72_wire(31 downto 0);
      type_cast_73_wire <= tmp_var; -- 
    end process;
    type_cast_91_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_91_inst_req_0;
      type_cast_91_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_91_inst_req_1;
      type_cast_91_inst_ack_1<= rack(0);
      type_cast_91_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_91_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_91_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_96_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_96_inst_req_0;
      type_cast_96_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_96_inst_req_1;
      type_cast_96_inst_ack_1<= rack(0);
      type_cast_96_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_96_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m2_factor_40,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_96_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_197_index_1_rename
    process(LSHR_u64_u64_196_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_196_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_196_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_index_1_resize
    process(LSHR_u64_u64_196_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_196_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_196_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_root_address_inst
    process(array_obj_ref_197_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_197_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_197_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_271_index_1_rename
    process(LSHR_u64_u64_270_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_270_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_270_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_271_index_1_resize
    process(LSHR_u64_u64_270_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_270_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_270_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_271_root_address_inst
    process(array_obj_ref_271_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_271_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_271_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_350_index_1_rename
    process(LSHR_u64_u64_349_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_349_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_349_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_350_index_1_resize
    process(LSHR_u64_u64_349_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_349_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_349_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_350_root_address_inst
    process(array_obj_ref_350_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_350_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_350_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_60_index_1_rename
    process(type_cast_59_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_59_resized;
      ov(13 downto 0) := iv;
      type_cast_59_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_60_index_1_resize
    process(type_cast_59_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_59_wire;
      ov := iv(13 downto 0);
      type_cast_59_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_60_root_address_inst
    process(array_obj_ref_60_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_60_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_60_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_74_index_1_rename
    process(type_cast_73_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_73_resized;
      ov(13 downto 0) := iv;
      type_cast_73_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_74_index_1_resize
    process(type_cast_73_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_73_wire;
      ov := iv(13 downto 0);
      type_cast_73_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_74_root_address_inst
    process(array_obj_ref_74_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_74_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_74_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_206_addr_0
    process(ptr_deref_206_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_206_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_206_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_206_base_resize
    process(fetch_addr1_199) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_199;
      ov := iv(13 downto 0);
      ptr_deref_206_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_206_gather_scatter
    process(ptr_deref_206_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_206_data_0;
      ov(63 downto 0) := iv;
      fv1_207 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_206_root_address_inst
    process(ptr_deref_206_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_206_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_206_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_280_addr_0
    process(ptr_deref_280_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_280_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_280_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_280_base_resize
    process(fetch_addr2_273) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_273;
      ov := iv(13 downto 0);
      ptr_deref_280_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_280_gather_scatter
    process(ptr_deref_280_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_280_data_0;
      ov(63 downto 0) := iv;
      fv2_281 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_280_root_address_inst
    process(ptr_deref_280_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_280_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_280_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_359_addr_0
    process(ptr_deref_359_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_359_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_359_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_359_base_resize
    process(fetch_addr3_352) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr3_352;
      ov := iv(13 downto 0);
      ptr_deref_359_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_359_gather_scatter
    process(ptr_deref_359_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_359_data_0;
      ov(63 downto 0) := iv;
      fv3_360 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_359_root_address_inst
    process(ptr_deref_359_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_359_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_359_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_51_addr_0
    process(ptr_deref_51_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_51_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_51_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_51_base_resize
    process(fetch_add1_48) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add1_48;
      ov := iv(13 downto 0);
      ptr_deref_51_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_51_gather_scatter
    process(ptr_deref_51_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_51_data_0;
      ov(63 downto 0) := iv;
      my_fetch1_52 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_51_root_address_inst
    process(ptr_deref_51_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_51_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_51_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_65_addr_0
    process(ptr_deref_65_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_65_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_65_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_65_base_resize
    process(fetch_add2_62) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add2_62;
      ov := iv(13 downto 0);
      ptr_deref_65_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_65_gather_scatter
    process(ptr_deref_65_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_65_data_0;
      ov(63 downto 0) := iv;
      my_fetch2_66 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_65_root_address_inst
    process(ptr_deref_65_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_65_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_65_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_79_addr_0
    process(ptr_deref_79_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_79_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_79_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_79_base_resize
    process(fetch_add3_76) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add3_76;
      ov := iv(13 downto 0);
      ptr_deref_79_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_79_gather_scatter
    process(ptr_deref_79_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_79_data_0;
      ov(63 downto 0) := iv;
      my_fetch3_80 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_79_root_address_inst
    process(ptr_deref_79_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_79_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_79_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_81_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_148;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_81_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_81_branch_req_0,
          ack0 => do_while_stmt_81_branch_ack_0,
          ack1 => do_while_stmt_81_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_168_inst
    process(row1_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row1_115, konst_167_wire_constant, tmp_var);
      ADD_u16_u16_168_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_242_inst
    process(row2_120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row2_120, konst_241_wire_constant, tmp_var);
      ADD_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_316_inst
    process(row3_125) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row3_125, konst_315_wire_constant, tmp_var);
      ADD_u16_u16_316_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_141_inst
    process(mycounter_98) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycounter_98, konst_140_wire_constant, tmp_var);
      ADD_u32_u32_141_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_175_inst
    process(address1_83) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_83, konst_174_wire_constant, tmp_var);
      n_address1_176 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_249_inst
    process(address2_88) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_88, konst_248_wire_constant, tmp_var);
      n_address2_250 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_323_inst
    process(address3_93) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address3_93, konst_322_wire_constant, tmp_var);
      n_address3_324 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_189_inst
    process(NEQ_u64_u1_187_wire, continue_185_delayed_1_0_179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_187_wire, continue_185_delayed_1_0_179, tmp_var);
      fn1_190 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_263_inst
    process(NEQ_u64_u1_261_wire, continue_247_delayed_1_0_253) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_261_wire, continue_247_delayed_1_0_253, tmp_var);
      fn2_264 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_337_inst
    process(NEQ_u64_u1_335_wire, continue_309_delayed_1_0_327) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_335_wire, continue_309_delayed_1_0_327, tmp_var);
      fn3_338 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_153_inst
    process(address1_83) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address1_83, konst_152_wire_constant, tmp_var);
      AND_u64_u64_153_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_227_inst
    process(address2_88) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address2_88, konst_226_wire_constant, tmp_var);
      AND_u64_u64_227_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_301_inst
    process(address3_93) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address3_93, konst_300_wire_constant, tmp_var);
      AND_u64_u64_301_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_134_inst
    process(mycounter_98, m_factor_35) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter_98, m_factor_35, tmp_var);
      next_row_135 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_58_inst
    process(m_factor_35) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_35, konst_57_wire_constant, tmp_var);
      LSHR_u32_u32_58_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_72_inst
    process(m_factor_35) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_35, konst_71_wire_constant, tmp_var);
      LSHR_u32_u32_72_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_161_inst
    process(fetch_val1_103, my_num1_157) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val1_103, my_num1_157, tmp_var);
      LSHR_u64_u64_161_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_183_inst
    process(n_address1_176) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_176, konst_182_wire_constant, tmp_var);
      LSHR_u64_u64_183_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_186_inst
    process(address1_83) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_83, konst_185_wire_constant, tmp_var);
      LSHR_u64_u64_186_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_196_inst
    process(n_address1_176) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_176, konst_195_wire_constant, tmp_var);
      LSHR_u64_u64_196_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_235_inst
    process(fetch_val2_107, my_num2_231) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val2_107, my_num2_231, tmp_var);
      LSHR_u64_u64_235_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_257_inst
    process(n_address2_250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_250, konst_256_wire_constant, tmp_var);
      LSHR_u64_u64_257_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_260_inst
    process(address2_88) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_88, konst_259_wire_constant, tmp_var);
      LSHR_u64_u64_260_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_270_inst
    process(n_address2_250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_250, konst_269_wire_constant, tmp_var);
      LSHR_u64_u64_270_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_309_inst
    process(fetch_val3_111, my_num3_305) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val3_111, my_num3_305, tmp_var);
      LSHR_u64_u64_309_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_331_inst
    process(n_address3_324) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_324, konst_330_wire_constant, tmp_var);
      LSHR_u64_u64_331_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_334_inst
    process(address3_93) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address3_93, konst_333_wire_constant, tmp_var);
      LSHR_u64_u64_334_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_349_inst
    process(n_address3_324) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_324, konst_348_wire_constant, tmp_var);
      LSHR_u64_u64_349_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_33_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_33_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_187_inst
    process(LSHR_u64_u64_183_wire, LSHR_u64_u64_186_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_183_wire, LSHR_u64_u64_186_wire, tmp_var);
      NEQ_u64_u1_187_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_261_inst
    process(LSHR_u64_u64_257_wire, LSHR_u64_u64_260_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_257_wire, LSHR_u64_u64_260_wire, tmp_var);
      NEQ_u64_u1_261_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_335_inst
    process(LSHR_u64_u64_331_wire, LSHR_u64_u64_334_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_331_wire, LSHR_u64_u64_334_wire, tmp_var);
      NEQ_u64_u1_335_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_39_inst
    process(m_factor_35) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(m_factor_35, konst_38_wire_constant, tmp_var);
      m2_factor_40 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_156_inst
    process(SUB_u64_u64_154_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_154_wire, konst_155_wire_constant, tmp_var);
      my_num1_157 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_230_inst
    process(SUB_u64_u64_228_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_228_wire, konst_229_wire_constant, tmp_var);
      my_num2_231 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_304_inst
    process(SUB_u64_u64_302_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_302_wire, konst_303_wire_constant, tmp_var);
      my_num3_305 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_154_inst
    process(konst_150_wire_constant, AND_u64_u64_153_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_150_wire_constant, AND_u64_u64_153_wire, tmp_var);
      SUB_u64_u64_154_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_228_inst
    process(konst_224_wire_constant, AND_u64_u64_227_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_224_wire_constant, AND_u64_u64_227_wire, tmp_var);
      SUB_u64_u64_228_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_302_inst
    process(konst_298_wire_constant, AND_u64_u64_301_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_298_wire_constant, AND_u64_u64_301_wire, tmp_var);
      SUB_u64_u64_302_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_147_inst
    process(n_row1_171, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row1_171, row_in_buffer, tmp_var);
      continue_148 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_342_inst
    process(row1_115, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row1_115, row_in_buffer, tmp_var);
      send_now3_343 <= tmp_var; --
    end process;
    -- shared split operator group (41) : array_obj_ref_197_index_offset 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_196_scaled;
      array_obj_ref_197_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_197_index_offset_req_0;
      array_obj_ref_197_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_197_index_offset_req_1;
      array_obj_ref_197_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_41_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_41_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : array_obj_ref_271_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_270_scaled;
      array_obj_ref_271_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_271_index_offset_req_0;
      array_obj_ref_271_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_271_index_offset_req_1;
      array_obj_ref_271_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : array_obj_ref_350_index_offset 
    ApIntAdd_group_43: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_349_scaled;
      array_obj_ref_350_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_350_index_offset_req_0;
      array_obj_ref_350_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_350_index_offset_req_1;
      array_obj_ref_350_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_43_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_43_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : array_obj_ref_60_index_offset 
    ApIntAdd_group_44: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_59_scaled;
      array_obj_ref_60_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_60_index_offset_req_0;
      array_obj_ref_60_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_60_index_offset_req_1;
      array_obj_ref_60_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_44_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : array_obj_ref_74_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_73_scaled;
      array_obj_ref_74_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_74_index_offset_req_0;
      array_obj_ref_74_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_74_index_offset_req_1;
      array_obj_ref_74_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared load operator group (0) : ptr_deref_79_load_0 ptr_deref_65_load_0 ptr_deref_206_load_0 ptr_deref_51_load_0 ptr_deref_280_load_0 ptr_deref_359_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(83 downto 0);
      signal data_out: std_logic_vector(383 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 2, 2 => 0, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 2, 2 => 1, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => true, 1 => true, 2 => false, 3 => true, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 6, 1 => 6, 2 => 2, 3 => 6, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_79_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_65_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_206_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_51_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_280_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_359_load_0_req_0;
      ptr_deref_79_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_65_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_206_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_51_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_280_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_359_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_79_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_65_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_206_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_51_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_280_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_359_load_0_req_1;
      ptr_deref_79_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_65_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_206_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_51_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_280_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_359_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn3_326_delayed_7_0_355(0);
      guard_vector(1)  <= fn2_259_delayed_7_0_276(0);
      guard_vector(2)  <=  '1';
      guard_vector(3)  <= fn1_197_delayed_7_0_202(0);
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 2) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_79_word_address_0 & ptr_deref_65_word_address_0 & ptr_deref_206_word_address_0 & ptr_deref_51_word_address_0 & ptr_deref_280_word_address_0 & ptr_deref_359_word_address_0;
      ptr_deref_79_data_0 <= data_out(383 downto 320);
      ptr_deref_65_data_0 <= data_out(319 downto 256);
      ptr_deref_206_data_0 <= data_out(255 downto 192);
      ptr_deref_51_data_0 <= data_out(191 downto 128);
      ptr_deref_280_data_0 <= data_out(127 downto 64);
      ptr_deref_359_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_220_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe1_220_inst_req_0;
      WPIPE_input_pipe1_220_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe1_220_inst_req_1;
      WPIPE_input_pipe1_220_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val1_163;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_input_pipe2_294_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe2_294_inst_req_0;
      WPIPE_input_pipe2_294_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe2_294_inst_req_1;
      WPIPE_input_pipe2_294_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val2_237;
      input_pipe2_write_1_gI: SplitGuardInterface generic map(name => "input_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "input_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe2_pipe_write_req(0),
          oack => input_pipe2_pipe_write_ack(0),
          odata => input_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_input_pipe3_374_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe3_374_inst_req_0;
      WPIPE_input_pipe3_374_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe3_374_inst_req_1;
      WPIPE_input_pipe3_374_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now3_343(0);
      data_in <= var_val3_311;
      input_pipe3_write_2_gI: SplitGuardInterface generic map(name => "input_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "input_pipe3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe3_pipe_write_req(0),
          oack => input_pipe3_pipe_write_ack(0),
          odata => input_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(47 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(63 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_3189_start: Boolean;
  signal convolution3D_CP_3189_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_1052_inst_ack_0 : boolean;
  signal type_cast_1056_inst_req_0 : boolean;
  signal type_cast_1056_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1052_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1052_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1065_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1065_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1077_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1065_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1065_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1115_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1115_inst_req_0 : boolean;
  signal type_cast_1119_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1090_inst_ack_0 : boolean;
  signal type_cast_1106_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1077_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1115_inst_ack_1 : boolean;
  signal type_cast_1106_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1090_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1115_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1102_inst_ack_1 : boolean;
  signal type_cast_1056_inst_req_1 : boolean;
  signal type_cast_1106_inst_ack_0 : boolean;
  signal type_cast_1056_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1090_inst_ack_1 : boolean;
  signal type_cast_1094_inst_ack_1 : boolean;
  signal type_cast_1094_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1077_inst_req_1 : boolean;
  signal type_cast_1081_inst_req_1 : boolean;
  signal type_cast_1069_inst_req_0 : boolean;
  signal type_cast_1069_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1102_inst_req_0 : boolean;
  signal type_cast_1094_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1102_inst_req_1 : boolean;
  signal type_cast_1481_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1052_inst_req_0 : boolean;
  signal type_cast_1081_inst_req_0 : boolean;
  signal type_cast_1106_inst_ack_1 : boolean;
  signal type_cast_1094_inst_ack_0 : boolean;
  signal type_cast_1081_inst_ack_1 : boolean;
  signal type_cast_1081_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1102_inst_ack_0 : boolean;
  signal type_cast_1069_inst_req_1 : boolean;
  signal type_cast_1069_inst_ack_1 : boolean;
  signal type_cast_1463_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1090_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1077_inst_req_0 : boolean;
  signal type_cast_1119_inst_ack_0 : boolean;
  signal type_cast_1119_inst_ack_1 : boolean;
  signal type_cast_1119_inst_req_1 : boolean;
  signal ptr_deref_1690_store_0_ack_0 : boolean;
  signal type_cast_1463_inst_req_1 : boolean;
  signal type_cast_1481_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2278_inst_ack_1 : boolean;
  signal type_cast_1782_inst_req_0 : boolean;
  signal type_cast_1782_inst_ack_0 : boolean;
  signal type_cast_1782_inst_req_1 : boolean;
  signal type_cast_1782_inst_ack_1 : boolean;
  signal type_cast_1705_inst_ack_1 : boolean;
  signal if_stmt_1572_branch_ack_0 : boolean;
  signal type_cast_2371_inst_ack_1 : boolean;
  signal type_cast_2371_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_2278_inst_req_1 : boolean;
  signal type_cast_2331_inst_ack_1 : boolean;
  signal type_cast_1791_inst_req_0 : boolean;
  signal type_cast_2299_inst_ack_1 : boolean;
  signal type_cast_1791_inst_ack_0 : boolean;
  signal type_cast_1773_inst_req_0 : boolean;
  signal type_cast_1764_inst_ack_0 : boolean;
  signal type_cast_1764_inst_req_1 : boolean;
  signal type_cast_1764_inst_ack_1 : boolean;
  signal type_cast_1773_inst_ack_0 : boolean;
  signal type_cast_1773_inst_req_1 : boolean;
  signal type_cast_1773_inst_ack_1 : boolean;
  signal type_cast_1463_inst_ack_1 : boolean;
  signal type_cast_1481_inst_req_1 : boolean;
  signal type_cast_1764_inst_req_0 : boolean;
  signal type_cast_1481_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_ack_1 : boolean;
  signal type_cast_1131_inst_req_0 : boolean;
  signal type_cast_1131_inst_ack_0 : boolean;
  signal type_cast_1131_inst_req_1 : boolean;
  signal type_cast_1131_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1140_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1140_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1140_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1140_inst_ack_1 : boolean;
  signal type_cast_1144_inst_req_0 : boolean;
  signal type_cast_1144_inst_ack_0 : boolean;
  signal type_cast_1144_inst_req_1 : boolean;
  signal type_cast_1144_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1152_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1152_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1152_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1152_inst_ack_1 : boolean;
  signal type_cast_1156_inst_req_0 : boolean;
  signal type_cast_1156_inst_ack_0 : boolean;
  signal type_cast_1156_inst_req_1 : boolean;
  signal type_cast_1156_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1165_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1165_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1165_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1165_inst_ack_1 : boolean;
  signal type_cast_1169_inst_req_0 : boolean;
  signal type_cast_1169_inst_ack_0 : boolean;
  signal type_cast_1169_inst_req_1 : boolean;
  signal type_cast_1169_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1177_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1177_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1177_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1177_inst_ack_1 : boolean;
  signal type_cast_1181_inst_req_0 : boolean;
  signal type_cast_1181_inst_ack_0 : boolean;
  signal type_cast_1181_inst_req_1 : boolean;
  signal type_cast_1181_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1190_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1190_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1190_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1190_inst_ack_1 : boolean;
  signal type_cast_1194_inst_req_0 : boolean;
  signal type_cast_1194_inst_ack_0 : boolean;
  signal type_cast_1194_inst_req_1 : boolean;
  signal type_cast_1194_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1202_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1202_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1202_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1202_inst_ack_1 : boolean;
  signal type_cast_1206_inst_req_0 : boolean;
  signal type_cast_1206_inst_ack_0 : boolean;
  signal type_cast_1206_inst_req_1 : boolean;
  signal type_cast_1206_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1215_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1215_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1215_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1215_inst_ack_1 : boolean;
  signal type_cast_1219_inst_req_0 : boolean;
  signal type_cast_1219_inst_ack_0 : boolean;
  signal type_cast_1219_inst_req_1 : boolean;
  signal type_cast_1219_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1227_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1227_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1227_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1227_inst_ack_1 : boolean;
  signal type_cast_1231_inst_req_0 : boolean;
  signal type_cast_1231_inst_ack_0 : boolean;
  signal type_cast_1231_inst_req_1 : boolean;
  signal if_stmt_1572_branch_ack_1 : boolean;
  signal type_cast_1231_inst_ack_1 : boolean;
  signal type_cast_1697_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1240_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1240_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1240_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1240_inst_ack_1 : boolean;
  signal type_cast_1705_inst_req_1 : boolean;
  signal type_cast_1701_inst_ack_0 : boolean;
  signal ptr_deref_1690_store_0_req_0 : boolean;
  signal type_cast_1640_inst_ack_1 : boolean;
  signal type_cast_1640_inst_req_1 : boolean;
  signal type_cast_1244_inst_req_0 : boolean;
  signal if_stmt_1572_branch_req_0 : boolean;
  signal type_cast_1244_inst_ack_0 : boolean;
  signal type_cast_1244_inst_req_1 : boolean;
  signal type_cast_1244_inst_ack_1 : boolean;
  signal type_cast_1697_inst_req_1 : boolean;
  signal if_stmt_1743_branch_ack_0 : boolean;
  signal WPIPE_num_out_pipe_2234_inst_req_1 : boolean;
  signal type_cast_1640_inst_ack_0 : boolean;
  signal type_cast_1640_inst_req_0 : boolean;
  signal type_cast_1253_inst_req_0 : boolean;
  signal type_cast_1253_inst_ack_0 : boolean;
  signal type_cast_1253_inst_req_1 : boolean;
  signal type_cast_1253_inst_ack_1 : boolean;
  signal type_cast_1697_inst_ack_0 : boolean;
  signal type_cast_1257_inst_req_0 : boolean;
  signal type_cast_1257_inst_ack_0 : boolean;
  signal type_cast_1257_inst_req_1 : boolean;
  signal type_cast_1257_inst_ack_1 : boolean;
  signal type_cast_1697_inst_req_0 : boolean;
  signal type_cast_1625_inst_ack_1 : boolean;
  signal type_cast_1625_inst_req_1 : boolean;
  signal type_cast_1272_inst_req_0 : boolean;
  signal type_cast_1272_inst_ack_0 : boolean;
  signal addr_of_1687_final_reg_ack_1 : boolean;
  signal type_cast_1272_inst_req_1 : boolean;
  signal if_stmt_1521_branch_ack_0 : boolean;
  signal type_cast_1272_inst_ack_1 : boolean;
  signal type_cast_1701_inst_ack_1 : boolean;
  signal if_stmt_1743_branch_ack_1 : boolean;
  signal type_cast_2401_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1477_inst_ack_1 : boolean;
  signal addr_of_1687_final_reg_req_1 : boolean;
  signal type_cast_1705_inst_ack_0 : boolean;
  signal type_cast_1463_inst_req_0 : boolean;
  signal if_stmt_1280_branch_req_0 : boolean;
  signal if_stmt_1280_branch_ack_1 : boolean;
  signal if_stmt_1280_branch_ack_0 : boolean;
  signal type_cast_1625_inst_ack_0 : boolean;
  signal type_cast_1300_inst_req_0 : boolean;
  signal type_cast_1300_inst_ack_0 : boolean;
  signal addr_of_1687_final_reg_ack_0 : boolean;
  signal addr_of_1687_final_reg_req_0 : boolean;
  signal type_cast_1300_inst_req_1 : boolean;
  signal type_cast_1300_inst_ack_1 : boolean;
  signal type_cast_1701_inst_req_1 : boolean;
  signal type_cast_1625_inst_req_0 : boolean;
  signal type_cast_1316_inst_req_0 : boolean;
  signal if_stmt_1521_branch_ack_1 : boolean;
  signal type_cast_1316_inst_ack_0 : boolean;
  signal type_cast_1316_inst_req_1 : boolean;
  signal type_cast_1316_inst_ack_1 : boolean;
  signal type_cast_1325_inst_req_0 : boolean;
  signal type_cast_1325_inst_ack_0 : boolean;
  signal type_cast_1325_inst_req_1 : boolean;
  signal if_stmt_1521_branch_req_0 : boolean;
  signal type_cast_1325_inst_ack_1 : boolean;
  signal if_stmt_1743_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_req_1 : boolean;
  signal type_cast_1335_inst_req_0 : boolean;
  signal type_cast_1335_inst_ack_0 : boolean;
  signal array_obj_ref_1686_index_offset_ack_1 : boolean;
  signal type_cast_1335_inst_req_1 : boolean;
  signal type_cast_1335_inst_ack_1 : boolean;
  signal ptr_deref_1690_store_0_ack_1 : boolean;
  signal ptr_deref_1690_store_0_req_1 : boolean;
  signal type_cast_2209_inst_ack_0 : boolean;
  signal if_stmt_1647_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_req_0 : boolean;
  signal type_cast_1701_inst_req_0 : boolean;
  signal type_cast_1499_inst_ack_1 : boolean;
  signal type_cast_1499_inst_req_1 : boolean;
  signal array_obj_ref_1370_index_offset_req_0 : boolean;
  signal array_obj_ref_1370_index_offset_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1477_inst_req_1 : boolean;
  signal array_obj_ref_1370_index_offset_req_1 : boolean;
  signal array_obj_ref_1370_index_offset_ack_1 : boolean;
  signal type_cast_1705_inst_req_0 : boolean;
  signal ptr_deref_1507_store_0_ack_1 : boolean;
  signal ptr_deref_1507_store_0_req_1 : boolean;
  signal array_obj_ref_1686_index_offset_req_1 : boolean;
  signal addr_of_1371_final_reg_req_0 : boolean;
  signal addr_of_1371_final_reg_ack_0 : boolean;
  signal addr_of_1371_final_reg_req_1 : boolean;
  signal addr_of_1371_final_reg_ack_1 : boolean;
  signal if_stmt_1647_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1374_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1374_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1374_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1374_inst_ack_1 : boolean;
  signal type_cast_1499_inst_ack_0 : boolean;
  signal type_cast_1499_inst_req_0 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal array_obj_ref_1686_index_offset_ack_0 : boolean;
  signal type_cast_1378_inst_req_1 : boolean;
  signal type_cast_1378_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1477_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1477_inst_req_0 : boolean;
  signal if_stmt_1647_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_req_0 : boolean;
  signal ptr_deref_1507_store_0_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_req_1 : boolean;
  signal ptr_deref_1507_store_0_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1495_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1495_inst_req_1 : boolean;
  signal array_obj_ref_1686_index_offset_req_0 : boolean;
  signal type_cast_1391_inst_req_0 : boolean;
  signal type_cast_1391_inst_ack_0 : boolean;
  signal type_cast_1391_inst_req_1 : boolean;
  signal type_cast_1391_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1495_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1495_inst_req_0 : boolean;
  signal type_cast_1409_inst_req_0 : boolean;
  signal type_cast_1409_inst_ack_0 : boolean;
  signal type_cast_1409_inst_req_1 : boolean;
  signal type_cast_1409_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2234_inst_ack_1 : boolean;
  signal call_stmt_2327_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1423_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1423_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1423_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1423_inst_ack_1 : boolean;
  signal type_cast_2351_inst_req_1 : boolean;
  signal type_cast_1427_inst_req_0 : boolean;
  signal type_cast_1427_inst_ack_0 : boolean;
  signal type_cast_1427_inst_req_1 : boolean;
  signal type_cast_1427_inst_ack_1 : boolean;
  signal type_cast_2199_inst_ack_1 : boolean;
  signal type_cast_2341_inst_req_0 : boolean;
  signal call_stmt_2327_call_ack_0 : boolean;
  signal call_stmt_2282_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1441_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1441_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1441_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1441_inst_ack_1 : boolean;
  signal type_cast_1445_inst_req_0 : boolean;
  signal type_cast_1445_inst_ack_0 : boolean;
  signal type_cast_1445_inst_req_1 : boolean;
  signal type_cast_1445_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_ack_1 : boolean;
  signal type_cast_1791_inst_req_1 : boolean;
  signal type_cast_1791_inst_ack_1 : boolean;
  signal type_cast_1796_inst_req_0 : boolean;
  signal type_cast_1796_inst_ack_0 : boolean;
  signal type_cast_1796_inst_req_1 : boolean;
  signal type_cast_1796_inst_ack_1 : boolean;
  signal type_cast_2209_inst_req_0 : boolean;
  signal type_cast_2299_inst_req_1 : boolean;
  signal array_obj_ref_1831_index_offset_req_0 : boolean;
  signal array_obj_ref_1831_index_offset_ack_0 : boolean;
  signal array_obj_ref_1831_index_offset_req_1 : boolean;
  signal array_obj_ref_1831_index_offset_ack_1 : boolean;
  signal call_stmt_2245_call_ack_0 : boolean;
  signal addr_of_1832_final_reg_req_0 : boolean;
  signal type_cast_2299_inst_ack_0 : boolean;
  signal addr_of_1832_final_reg_ack_0 : boolean;
  signal call_stmt_2245_call_req_0 : boolean;
  signal type_cast_2371_inst_ack_0 : boolean;
  signal addr_of_1832_final_reg_req_1 : boolean;
  signal type_cast_2299_inst_req_0 : boolean;
  signal addr_of_1832_final_reg_ack_1 : boolean;
  signal type_cast_2401_inst_req_0 : boolean;
  signal type_cast_2331_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_2278_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2278_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1835_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1835_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1835_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1835_inst_ack_1 : boolean;
  signal type_cast_2391_inst_ack_1 : boolean;
  signal type_cast_2391_inst_req_1 : boolean;
  signal type_cast_2351_inst_ack_1 : boolean;
  signal type_cast_2371_inst_req_0 : boolean;
  signal type_cast_1839_inst_req_0 : boolean;
  signal type_cast_1839_inst_ack_0 : boolean;
  signal type_cast_1839_inst_req_1 : boolean;
  signal type_cast_1839_inst_ack_1 : boolean;
  signal type_cast_2401_inst_req_1 : boolean;
  signal type_cast_2331_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1848_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1848_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_2234_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1848_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1848_inst_ack_1 : boolean;
  signal type_cast_2391_inst_ack_0 : boolean;
  signal type_cast_2391_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_2274_inst_ack_1 : boolean;
  signal type_cast_1852_inst_req_0 : boolean;
  signal type_cast_2295_inst_ack_1 : boolean;
  signal type_cast_1852_inst_ack_0 : boolean;
  signal type_cast_1852_inst_req_1 : boolean;
  signal type_cast_2295_inst_req_1 : boolean;
  signal type_cast_1852_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2234_inst_req_0 : boolean;
  signal type_cast_2331_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_2274_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1866_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1866_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1866_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1866_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_2274_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2274_inst_req_0 : boolean;
  signal type_cast_2295_inst_ack_0 : boolean;
  signal type_cast_1870_inst_req_0 : boolean;
  signal type_cast_1870_inst_ack_0 : boolean;
  signal type_cast_2295_inst_req_0 : boolean;
  signal type_cast_1870_inst_req_1 : boolean;
  signal type_cast_1870_inst_ack_1 : boolean;
  signal type_cast_2351_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1884_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1884_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1884_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1884_inst_ack_1 : boolean;
  signal type_cast_2271_inst_ack_1 : boolean;
  signal type_cast_2271_inst_req_1 : boolean;
  signal type_cast_1888_inst_req_0 : boolean;
  signal type_cast_1888_inst_ack_0 : boolean;
  signal type_cast_1888_inst_req_1 : boolean;
  signal type_cast_2199_inst_req_1 : boolean;
  signal type_cast_1888_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2231_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2231_inst_req_1 : boolean;
  signal type_cast_2351_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1902_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1902_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1902_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1902_inst_ack_1 : boolean;
  signal type_cast_2271_inst_ack_0 : boolean;
  signal type_cast_2381_inst_ack_1 : boolean;
  signal type_cast_2381_inst_req_1 : boolean;
  signal type_cast_2271_inst_req_0 : boolean;
  signal type_cast_1906_inst_req_0 : boolean;
  signal type_cast_1906_inst_ack_0 : boolean;
  signal type_cast_1906_inst_req_1 : boolean;
  signal type_cast_2286_inst_ack_1 : boolean;
  signal type_cast_1906_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2231_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1920_inst_req_0 : boolean;
  signal type_cast_2286_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1920_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_2231_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1920_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1920_inst_ack_1 : boolean;
  signal if_stmt_2261_branch_ack_0 : boolean;
  signal type_cast_2361_inst_ack_1 : boolean;
  signal type_cast_1924_inst_req_0 : boolean;
  signal type_cast_1924_inst_ack_0 : boolean;
  signal type_cast_2361_inst_req_1 : boolean;
  signal type_cast_1924_inst_req_1 : boolean;
  signal type_cast_2286_inst_ack_0 : boolean;
  signal type_cast_1924_inst_ack_1 : boolean;
  signal type_cast_2341_inst_ack_1 : boolean;
  signal type_cast_2341_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1938_inst_req_0 : boolean;
  signal type_cast_2286_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1938_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1938_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1938_inst_ack_1 : boolean;
  signal type_cast_2381_inst_ack_0 : boolean;
  signal if_stmt_2261_branch_ack_1 : boolean;
  signal type_cast_1942_inst_req_0 : boolean;
  signal type_cast_1942_inst_ack_0 : boolean;
  signal type_cast_1942_inst_req_1 : boolean;
  signal type_cast_1942_inst_ack_1 : boolean;
  signal call_stmt_2327_call_ack_1 : boolean;
  signal call_stmt_2327_call_req_1 : boolean;
  signal type_cast_2341_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1956_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1956_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1956_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1956_inst_ack_1 : boolean;
  signal if_stmt_2261_branch_req_0 : boolean;
  signal type_cast_2381_inst_req_0 : boolean;
  signal type_cast_2361_inst_ack_0 : boolean;
  signal type_cast_1960_inst_req_0 : boolean;
  signal type_cast_1960_inst_ack_0 : boolean;
  signal type_cast_2361_inst_req_0 : boolean;
  signal type_cast_1960_inst_req_1 : boolean;
  signal call_stmt_2282_call_ack_1 : boolean;
  signal type_cast_1960_inst_ack_1 : boolean;
  signal type_cast_2209_inst_ack_1 : boolean;
  signal call_stmt_2249_call_ack_1 : boolean;
  signal call_stmt_2249_call_req_1 : boolean;
  signal call_stmt_2249_call_ack_0 : boolean;
  signal call_stmt_2249_call_req_0 : boolean;
  signal call_stmt_2282_call_req_1 : boolean;
  signal type_cast_2209_inst_req_1 : boolean;
  signal call_stmt_2282_call_ack_0 : boolean;
  signal ptr_deref_1968_store_0_req_0 : boolean;
  signal call_stmt_2245_call_ack_1 : boolean;
  signal ptr_deref_1968_store_0_ack_0 : boolean;
  signal ptr_deref_1968_store_0_req_1 : boolean;
  signal call_stmt_2245_call_req_1 : boolean;
  signal ptr_deref_1968_store_0_ack_1 : boolean;
  signal if_stmt_1982_branch_req_0 : boolean;
  signal if_stmt_1982_branch_ack_1 : boolean;
  signal if_stmt_1982_branch_ack_0 : boolean;
  signal if_stmt_2033_branch_req_0 : boolean;
  signal if_stmt_2033_branch_ack_1 : boolean;
  signal if_stmt_2033_branch_ack_0 : boolean;
  signal type_cast_2048_inst_req_0 : boolean;
  signal type_cast_2048_inst_ack_0 : boolean;
  signal type_cast_2048_inst_req_1 : boolean;
  signal type_cast_2048_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2086_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2086_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2086_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2086_inst_ack_1 : boolean;
  signal type_cast_2090_inst_req_0 : boolean;
  signal type_cast_2090_inst_ack_0 : boolean;
  signal type_cast_2090_inst_req_1 : boolean;
  signal type_cast_2090_inst_ack_1 : boolean;
  signal type_cast_2105_inst_req_0 : boolean;
  signal type_cast_2105_inst_ack_0 : boolean;
  signal type_cast_2105_inst_req_1 : boolean;
  signal type_cast_2105_inst_ack_1 : boolean;
  signal if_stmt_2112_branch_req_0 : boolean;
  signal if_stmt_2112_branch_ack_1 : boolean;
  signal if_stmt_2112_branch_ack_0 : boolean;
  signal array_obj_ref_2151_index_offset_req_0 : boolean;
  signal array_obj_ref_2151_index_offset_ack_0 : boolean;
  signal array_obj_ref_2151_index_offset_req_1 : boolean;
  signal array_obj_ref_2151_index_offset_ack_1 : boolean;
  signal addr_of_2152_final_reg_req_0 : boolean;
  signal addr_of_2152_final_reg_ack_0 : boolean;
  signal addr_of_2152_final_reg_req_1 : boolean;
  signal addr_of_2152_final_reg_ack_1 : boolean;
  signal ptr_deref_2155_store_0_req_0 : boolean;
  signal ptr_deref_2155_store_0_ack_0 : boolean;
  signal ptr_deref_2155_store_0_req_1 : boolean;
  signal ptr_deref_2155_store_0_ack_1 : boolean;
  signal ptr_deref_2169_store_0_req_0 : boolean;
  signal ptr_deref_2169_store_0_ack_0 : boolean;
  signal ptr_deref_2169_store_0_req_1 : boolean;
  signal ptr_deref_2169_store_0_ack_1 : boolean;
  signal call_stmt_2175_call_req_0 : boolean;
  signal call_stmt_2175_call_ack_0 : boolean;
  signal call_stmt_2175_call_req_1 : boolean;
  signal call_stmt_2175_call_ack_1 : boolean;
  signal WPIPE_output_pipe_2176_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2176_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_2176_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2176_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2179_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2179_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_2179_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2179_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2182_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2182_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_2182_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2182_inst_ack_1 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal type_cast_2401_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2403_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2403_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2403_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2403_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2406_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2406_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2406_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2406_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2409_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2409_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2409_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2409_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2412_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2412_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2412_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2412_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2415_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2415_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2415_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2415_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2418_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2418_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2418_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2418_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2421_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2421_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2421_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2421_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2424_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2424_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2424_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2424_inst_ack_1 : boolean;
  signal phi_stmt_1358_req_0 : boolean;
  signal type_cast_1364_inst_req_0 : boolean;
  signal type_cast_1364_inst_ack_0 : boolean;
  signal type_cast_1364_inst_req_1 : boolean;
  signal type_cast_1364_inst_ack_1 : boolean;
  signal phi_stmt_1358_req_1 : boolean;
  signal phi_stmt_1358_ack_0 : boolean;
  signal phi_stmt_1552_req_1 : boolean;
  signal type_cast_1555_inst_req_0 : boolean;
  signal type_cast_1555_inst_ack_0 : boolean;
  signal type_cast_1555_inst_req_1 : boolean;
  signal type_cast_1555_inst_ack_1 : boolean;
  signal phi_stmt_1552_req_0 : boolean;
  signal phi_stmt_1552_ack_0 : boolean;
  signal phi_stmt_1593_req_0 : boolean;
  signal phi_stmt_1600_req_0 : boolean;
  signal type_cast_1599_inst_req_0 : boolean;
  signal type_cast_1599_inst_ack_0 : boolean;
  signal type_cast_1599_inst_req_1 : boolean;
  signal type_cast_1599_inst_ack_1 : boolean;
  signal phi_stmt_1593_req_1 : boolean;
  signal type_cast_1606_inst_req_0 : boolean;
  signal type_cast_1606_inst_ack_0 : boolean;
  signal type_cast_1606_inst_req_1 : boolean;
  signal type_cast_1606_inst_ack_1 : boolean;
  signal phi_stmt_1600_req_1 : boolean;
  signal phi_stmt_1593_ack_0 : boolean;
  signal phi_stmt_1600_ack_0 : boolean;
  signal type_cast_1657_inst_req_0 : boolean;
  signal type_cast_1657_inst_ack_0 : boolean;
  signal type_cast_1657_inst_req_1 : boolean;
  signal type_cast_1657_inst_ack_1 : boolean;
  signal phi_stmt_1654_req_0 : boolean;
  signal phi_stmt_1654_ack_0 : boolean;
  signal phi_stmt_1819_req_1 : boolean;
  signal type_cast_1822_inst_req_0 : boolean;
  signal type_cast_1822_inst_ack_0 : boolean;
  signal type_cast_1822_inst_req_1 : boolean;
  signal type_cast_1822_inst_ack_1 : boolean;
  signal phi_stmt_1819_req_0 : boolean;
  signal phi_stmt_1819_ack_0 : boolean;
  signal type_cast_2016_inst_req_0 : boolean;
  signal type_cast_2016_inst_ack_0 : boolean;
  signal type_cast_2016_inst_req_1 : boolean;
  signal type_cast_2016_inst_ack_1 : boolean;
  signal phi_stmt_2013_req_0 : boolean;
  signal phi_stmt_2013_req_1 : boolean;
  signal phi_stmt_2013_ack_0 : boolean;
  signal phi_stmt_2065_req_1 : boolean;
  signal phi_stmt_2058_req_1 : boolean;
  signal type_cast_2068_inst_req_0 : boolean;
  signal type_cast_2068_inst_ack_0 : boolean;
  signal type_cast_2068_inst_req_1 : boolean;
  signal type_cast_2068_inst_ack_1 : boolean;
  signal phi_stmt_2065_req_0 : boolean;
  signal type_cast_2061_inst_req_0 : boolean;
  signal type_cast_2061_inst_ack_0 : boolean;
  signal type_cast_2061_inst_req_1 : boolean;
  signal type_cast_2061_inst_ack_1 : boolean;
  signal phi_stmt_2058_req_0 : boolean;
  signal phi_stmt_2058_ack_0 : boolean;
  signal phi_stmt_2065_ack_0 : boolean;
  signal type_cast_2122_inst_req_0 : boolean;
  signal type_cast_2122_inst_ack_0 : boolean;
  signal type_cast_2122_inst_req_1 : boolean;
  signal type_cast_2122_inst_ack_1 : boolean;
  signal phi_stmt_2119_req_0 : boolean;
  signal phi_stmt_2119_ack_0 : boolean;
  signal phi_stmt_2218_req_0 : boolean;
  signal type_cast_2224_inst_req_0 : boolean;
  signal type_cast_2224_inst_ack_0 : boolean;
  signal type_cast_2224_inst_req_1 : boolean;
  signal type_cast_2224_inst_ack_1 : boolean;
  signal phi_stmt_2218_req_1 : boolean;
  signal phi_stmt_2218_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_3189_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3189_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_3189_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3189_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_3189: Block -- control-path 
    signal convolution3D_CP_3189_elements: BooleanArray(382 downto 0);
    -- 
  begin -- 
    convolution3D_CP_3189_elements(0) <= convolution3D_CP_3189_start;
    convolution3D_CP_3189_symbol <= convolution3D_CP_3189_elements(313);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1049/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/branch_block_stmt_1049__entry__
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279__entry__
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Update/cr
      -- 
    cr_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1106_inst_req_1); -- 
    cr_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1056_inst_req_1); -- 
    cr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1094_inst_req_1); -- 
    cr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1081_inst_req_1); -- 
    rr_3311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => RPIPE_maxpool_input_pipe_1052_inst_req_0); -- 
    cr_3358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1069_inst_req_1); -- 
    cr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1119_inst_req_1); -- 
    cr_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1131_inst_req_1); -- 
    cr_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1144_inst_req_1); -- 
    cr_3554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1156_inst_req_1); -- 
    cr_3582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1169_inst_req_1); -- 
    cr_3610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1181_inst_req_1); -- 
    cr_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1194_inst_req_1); -- 
    cr_3666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1206_inst_req_1); -- 
    cr_3694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1219_inst_req_1); -- 
    cr_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1231_inst_req_1); -- 
    cr_3750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1244_inst_req_1); -- 
    cr_3764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1253_inst_req_1); -- 
    cr_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1257_inst_req_1); -- 
    cr_3792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(0), ack => type_cast_1272_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Sample/$exit
      -- 
    ra_3312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1052_inst_ack_0, ack => convolution3D_CP_3189_elements(1)); -- 
    cr_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(1), ack => RPIPE_maxpool_input_pipe_1052_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1052_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_sample_start_
      -- 
    ca_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1052_inst_ack_1, ack => convolution3D_CP_3189_elements(2)); -- 
    rr_3325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(2), ack => type_cast_1056_inst_req_0); -- 
    rr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(2), ack => RPIPE_maxpool_input_pipe_1065_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Sample/$exit
      -- 
    ra_3326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_0, ack => convolution3D_CP_3189_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1056_Update/ca
      -- 
    ca_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_1, ack => convolution3D_CP_3189_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_update_start_
      -- 
    ra_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1065_inst_ack_0, ack => convolution3D_CP_3189_elements(5)); -- 
    cr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(5), ack => RPIPE_maxpool_input_pipe_1065_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1065_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Sample/rr
      -- 
    ca_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1065_inst_ack_1, ack => convolution3D_CP_3189_elements(6)); -- 
    rr_3353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(6), ack => type_cast_1069_inst_req_0); -- 
    rr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(6), ack => RPIPE_maxpool_input_pipe_1077_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Sample/ra
      -- 
    ra_3354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1069_inst_ack_0, ack => convolution3D_CP_3189_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1069_Update/ca
      -- 
    ca_3359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1069_inst_ack_1, ack => convolution3D_CP_3189_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Sample/$exit
      -- 
    ra_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1077_inst_ack_0, ack => convolution3D_CP_3189_elements(9)); -- 
    cr_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(9), ack => RPIPE_maxpool_input_pipe_1077_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1077_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Sample/rr
      -- 
    ca_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1077_inst_ack_1, ack => convolution3D_CP_3189_elements(10)); -- 
    rr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(10), ack => type_cast_1081_inst_req_0); -- 
    rr_3395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(10), ack => RPIPE_maxpool_input_pipe_1090_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Sample/ra
      -- 
    ra_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1081_inst_ack_0, ack => convolution3D_CP_3189_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1081_Update/ca
      -- 
    ca_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1081_inst_ack_1, ack => convolution3D_CP_3189_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_update_start_
      -- 
    ra_3396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1090_inst_ack_0, ack => convolution3D_CP_3189_elements(13)); -- 
    cr_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(13), ack => RPIPE_maxpool_input_pipe_1090_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1090_Update/$exit
      -- 
    ca_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1090_inst_ack_1, ack => convolution3D_CP_3189_elements(14)); -- 
    rr_3423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(14), ack => RPIPE_maxpool_input_pipe_1102_inst_req_0); -- 
    rr_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(14), ack => type_cast_1094_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Sample/ra
      -- 
    ra_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1094_inst_ack_0, ack => convolution3D_CP_3189_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1094_update_completed_
      -- 
    ca_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1094_inst_ack_1, ack => convolution3D_CP_3189_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_update_start_
      -- 
    ra_3424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1102_inst_ack_0, ack => convolution3D_CP_3189_elements(17)); -- 
    cr_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(17), ack => RPIPE_maxpool_input_pipe_1102_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1102_update_completed_
      -- 
    ca_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1102_inst_ack_1, ack => convolution3D_CP_3189_elements(18)); -- 
    rr_3451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(18), ack => RPIPE_maxpool_input_pipe_1115_inst_req_0); -- 
    rr_3437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(18), ack => type_cast_1106_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_sample_completed_
      -- 
    ra_3438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_0, ack => convolution3D_CP_3189_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1106_update_completed_
      -- 
    ca_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_1, ack => convolution3D_CP_3189_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_update_start_
      -- 
    ra_3452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1115_inst_ack_0, ack => convolution3D_CP_3189_elements(21)); -- 
    cr_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(21), ack => RPIPE_maxpool_input_pipe_1115_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1115_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Sample/rr
      -- 
    ca_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1115_inst_ack_1, ack => convolution3D_CP_3189_elements(22)); -- 
    rr_3479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(22), ack => RPIPE_maxpool_input_pipe_1127_inst_req_0); -- 
    rr_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(22), ack => type_cast_1119_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Sample/ra
      -- 
    ra_3466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1119_inst_ack_0, ack => convolution3D_CP_3189_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1119_Update/$exit
      -- 
    ca_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1119_inst_ack_1, ack => convolution3D_CP_3189_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Update/cr
      -- 
    ra_3480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1127_inst_ack_0, ack => convolution3D_CP_3189_elements(25)); -- 
    cr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(25), ack => RPIPE_maxpool_input_pipe_1127_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1127_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Sample/rr
      -- 
    ca_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1127_inst_ack_1, ack => convolution3D_CP_3189_elements(26)); -- 
    rr_3493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(26), ack => type_cast_1131_inst_req_0); -- 
    rr_3507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(26), ack => RPIPE_maxpool_input_pipe_1140_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Sample/ra
      -- 
    ra_3494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_0, ack => convolution3D_CP_3189_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1131_Update/ca
      -- 
    ca_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_1, ack => convolution3D_CP_3189_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Update/cr
      -- 
    ra_3508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1140_inst_ack_0, ack => convolution3D_CP_3189_elements(29)); -- 
    cr_3512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(29), ack => RPIPE_maxpool_input_pipe_1140_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1140_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Sample/rr
      -- 
    ca_3513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1140_inst_ack_1, ack => convolution3D_CP_3189_elements(30)); -- 
    rr_3521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(30), ack => type_cast_1144_inst_req_0); -- 
    rr_3535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(30), ack => RPIPE_maxpool_input_pipe_1152_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Sample/ra
      -- 
    ra_3522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1144_inst_ack_0, ack => convolution3D_CP_3189_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1144_Update/ca
      -- 
    ca_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1144_inst_ack_1, ack => convolution3D_CP_3189_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Update/cr
      -- 
    ra_3536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1152_inst_ack_0, ack => convolution3D_CP_3189_elements(33)); -- 
    cr_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(33), ack => RPIPE_maxpool_input_pipe_1152_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1152_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Sample/rr
      -- 
    ca_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1152_inst_ack_1, ack => convolution3D_CP_3189_elements(34)); -- 
    rr_3549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(34), ack => type_cast_1156_inst_req_0); -- 
    rr_3563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(34), ack => RPIPE_maxpool_input_pipe_1165_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Sample/ra
      -- 
    ra_3550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_0, ack => convolution3D_CP_3189_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1156_Update/ca
      -- 
    ca_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_1, ack => convolution3D_CP_3189_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Update/cr
      -- 
    ra_3564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1165_inst_ack_0, ack => convolution3D_CP_3189_elements(37)); -- 
    cr_3568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(37), ack => RPIPE_maxpool_input_pipe_1165_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1165_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Sample/rr
      -- 
    ca_3569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1165_inst_ack_1, ack => convolution3D_CP_3189_elements(38)); -- 
    rr_3591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(38), ack => RPIPE_maxpool_input_pipe_1177_inst_req_0); -- 
    rr_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(38), ack => type_cast_1169_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Sample/ra
      -- 
    ra_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_0, ack => convolution3D_CP_3189_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1169_Update/ca
      -- 
    ca_3583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_1, ack => convolution3D_CP_3189_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Update/cr
      -- 
    ra_3592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1177_inst_ack_0, ack => convolution3D_CP_3189_elements(41)); -- 
    cr_3596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(41), ack => RPIPE_maxpool_input_pipe_1177_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1177_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Sample/rr
      -- 
    ca_3597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1177_inst_ack_1, ack => convolution3D_CP_3189_elements(42)); -- 
    rr_3605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(42), ack => type_cast_1181_inst_req_0); -- 
    rr_3619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(42), ack => RPIPE_maxpool_input_pipe_1190_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Sample/ra
      -- 
    ra_3606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1181_inst_ack_0, ack => convolution3D_CP_3189_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1181_Update/ca
      -- 
    ca_3611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1181_inst_ack_1, ack => convolution3D_CP_3189_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Update/cr
      -- 
    ra_3620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1190_inst_ack_0, ack => convolution3D_CP_3189_elements(45)); -- 
    cr_3624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(45), ack => RPIPE_maxpool_input_pipe_1190_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1190_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Sample/rr
      -- 
    ca_3625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1190_inst_ack_1, ack => convolution3D_CP_3189_elements(46)); -- 
    rr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(46), ack => RPIPE_maxpool_input_pipe_1202_inst_req_0); -- 
    rr_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(46), ack => type_cast_1194_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Sample/ra
      -- 
    ra_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1194_inst_ack_0, ack => convolution3D_CP_3189_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1194_Update/ca
      -- 
    ca_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1194_inst_ack_1, ack => convolution3D_CP_3189_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Update/cr
      -- 
    ra_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1202_inst_ack_0, ack => convolution3D_CP_3189_elements(49)); -- 
    cr_3652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(49), ack => RPIPE_maxpool_input_pipe_1202_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1202_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Sample/rr
      -- 
    ca_3653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1202_inst_ack_1, ack => convolution3D_CP_3189_elements(50)); -- 
    rr_3661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(50), ack => type_cast_1206_inst_req_0); -- 
    rr_3675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(50), ack => RPIPE_maxpool_input_pipe_1215_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Sample/ra
      -- 
    ra_3662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_0, ack => convolution3D_CP_3189_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1206_Update/ca
      -- 
    ca_3667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_1, ack => convolution3D_CP_3189_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Update/cr
      -- 
    ra_3676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1215_inst_ack_0, ack => convolution3D_CP_3189_elements(53)); -- 
    cr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(53), ack => RPIPE_maxpool_input_pipe_1215_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1215_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Sample/rr
      -- 
    ca_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1215_inst_ack_1, ack => convolution3D_CP_3189_elements(54)); -- 
    rr_3689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(54), ack => type_cast_1219_inst_req_0); -- 
    rr_3703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(54), ack => RPIPE_maxpool_input_pipe_1227_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Sample/ra
      -- 
    ra_3690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_0, ack => convolution3D_CP_3189_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1219_Update/ca
      -- 
    ca_3695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_1, ack => convolution3D_CP_3189_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Update/cr
      -- 
    ra_3704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1227_inst_ack_0, ack => convolution3D_CP_3189_elements(57)); -- 
    cr_3708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(57), ack => RPIPE_maxpool_input_pipe_1227_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1227_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Sample/rr
      -- 
    ca_3709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1227_inst_ack_1, ack => convolution3D_CP_3189_elements(58)); -- 
    rr_3717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(58), ack => type_cast_1231_inst_req_0); -- 
    rr_3731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(58), ack => RPIPE_maxpool_input_pipe_1240_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Sample/ra
      -- 
    ra_3718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_0, ack => convolution3D_CP_3189_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1231_Update/ca
      -- 
    ca_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_1, ack => convolution3D_CP_3189_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_update_start_
      -- CP-element group 61: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Update/cr
      -- 
    ra_3732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1240_inst_ack_0, ack => convolution3D_CP_3189_elements(61)); -- 
    cr_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(61), ack => RPIPE_maxpool_input_pipe_1240_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/RPIPE_maxpool_input_pipe_1240_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Sample/rr
      -- 
    ca_3737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1240_inst_ack_1, ack => convolution3D_CP_3189_elements(62)); -- 
    rr_3745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(62), ack => type_cast_1244_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Sample/ra
      -- 
    ra_3746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1244_inst_ack_0, ack => convolution3D_CP_3189_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1244_Update/ca
      -- 
    ca_3751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1244_inst_ack_1, ack => convolution3D_CP_3189_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	16 
    -- CP-element group 65: 	12 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Sample/rr
      -- 
    rr_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(65), ack => type_cast_1253_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(16) & convolution3D_CP_3189_elements(12);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Sample/ra
      -- 
    ra_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_0, ack => convolution3D_CP_3189_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1253_Update/ca
      -- 
    ca_3765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_1, ack => convolution3D_CP_3189_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Sample/rr
      -- 
    rr_3773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(68), ack => type_cast_1257_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(20) & convolution3D_CP_3189_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Sample/ra
      -- 
    ra_3774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1257_inst_ack_0, ack => convolution3D_CP_3189_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1257_Update/ca
      -- 
    ca_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1257_inst_ack_1, ack => convolution3D_CP_3189_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Sample/rr
      -- 
    rr_3787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(71), ack => type_cast_1272_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(67) & convolution3D_CP_3189_elements(70) & convolution3D_CP_3189_elements(4) & convolution3D_CP_3189_elements(8);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Sample/ra
      -- 
    ra_3788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1272_inst_ack_0, ack => convolution3D_CP_3189_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/type_cast_1272_Update/ca
      -- 
    ca_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1272_inst_ack_1, ack => convolution3D_CP_3189_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	28 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279/$exit
      -- CP-element group 74: 	 branch_block_stmt_1049/assign_stmt_1053_to_assign_stmt_1279__exit__
      -- CP-element group 74: 	 branch_block_stmt_1049/if_stmt_1280__entry__
      -- CP-element group 74: 	 branch_block_stmt_1049/if_stmt_1280_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1049/if_stmt_1280_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1049/if_stmt_1280_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1049/if_stmt_1280_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1049/R_cmp383_1281_place
      -- CP-element group 74: 	 branch_block_stmt_1049/if_stmt_1280_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1049/if_stmt_1280_else_link/$entry
      -- 
    branch_req_3801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(74), ack => if_stmt_1280_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(40) & convolution3D_CP_3189_elements(32) & convolution3D_CP_3189_elements(36) & convolution3D_CP_3189_elements(44) & convolution3D_CP_3189_elements(48) & convolution3D_CP_3189_elements(52) & convolution3D_CP_3189_elements(56) & convolution3D_CP_3189_elements(60) & convolution3D_CP_3189_elements(64) & convolution3D_CP_3189_elements(73) & convolution3D_CP_3189_elements(28);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_1049/merge_stmt_1286__exit__
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355__entry__
      -- CP-element group 75: 	 branch_block_stmt_1049/if_stmt_1280_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1049/if_stmt_1280_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1049/entry_bbx_xnph385
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1049/entry_bbx_xnph385_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/entry_bbx_xnph385_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1049/merge_stmt_1286_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1049/merge_stmt_1286_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1049/merge_stmt_1286_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1049/merge_stmt_1286_PhiAck/dummy
      -- 
    if_choice_transition_3806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1280_branch_ack_1, ack => convolution3D_CP_3189_elements(75)); -- 
    rr_3823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(75), ack => type_cast_1300_inst_req_0); -- 
    cr_3828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(75), ack => type_cast_1300_inst_req_1); -- 
    rr_3837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(75), ack => type_cast_1316_inst_req_0); -- 
    cr_3842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(75), ack => type_cast_1316_inst_req_1); -- 
    rr_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(75), ack => type_cast_1325_inst_req_0); -- 
    cr_3856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(75), ack => type_cast_1325_inst_req_1); -- 
    cr_3870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(75), ack => type_cast_1335_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	320 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_1049/if_stmt_1280_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1049/if_stmt_1280_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1049/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/phi_stmt_1552/$entry
      -- CP-element group 76: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$entry
      -- 
    else_choice_transition_3810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1280_branch_ack_0, ack => convolution3D_CP_3189_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Sample/ra
      -- 
    ra_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_0, ack => convolution3D_CP_3189_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1300_Update/ca
      -- 
    ca_3829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_1, ack => convolution3D_CP_3189_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Sample/ra
      -- 
    ra_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_0, ack => convolution3D_CP_3189_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1316_Update/ca
      -- 
    ca_3843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_1, ack => convolution3D_CP_3189_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Sample/ra
      -- 
    ra_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_0, ack => convolution3D_CP_3189_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1325_Update/ca
      -- 
    ca_3857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_1, ack => convolution3D_CP_3189_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Sample/rr
      -- 
    rr_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(83), ack => type_cast_1335_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(80) & convolution3D_CP_3189_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Sample/ra
      -- 
    ra_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1335_inst_ack_0, ack => convolution3D_CP_3189_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/type_cast_1335_Update/ca
      -- 
    ca_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1335_inst_ack_1, ack => convolution3D_CP_3189_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	314 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355__exit__
      -- CP-element group 86: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_1049/assign_stmt_1291_to_assign_stmt_1355/$exit
      -- CP-element group 86: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1358/$entry
      -- CP-element group 86: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(78) & convolution3D_CP_3189_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	319 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Sample/ack
      -- 
    ack_3900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1370_index_offset_ack_0, ack => convolution3D_CP_3189_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	319 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_request/req
      -- 
    ack_3905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1370_index_offset_ack_1, ack => convolution3D_CP_3189_elements(88)); -- 
    req_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(88), ack => addr_of_1371_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_request/ack
      -- 
    ack_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1371_final_reg_ack_0, ack => convolution3D_CP_3189_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	319 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_word_addrgen/root_register_ack
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_complete/ack
      -- 
    ack_3920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1371_final_reg_ack_1, ack => convolution3D_CP_3189_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	319 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Update/cr
      -- 
    ra_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1374_inst_ack_0, ack => convolution3D_CP_3189_elements(91)); -- 
    cr_3933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(91), ack => RPIPE_maxpool_input_pipe_1374_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Sample/rr
      -- 
    ca_3934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1374_inst_ack_1, ack => convolution3D_CP_3189_elements(92)); -- 
    rr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(92), ack => type_cast_1378_inst_req_0); -- 
    rr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(92), ack => RPIPE_maxpool_input_pipe_1387_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Sample/ra
      -- 
    ra_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_0, ack => convolution3D_CP_3189_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	319 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Update/ca
      -- 
    ca_3948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_1, ack => convolution3D_CP_3189_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_update_start_
      -- CP-element group 95: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Update/cr
      -- 
    ra_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1387_inst_ack_0, ack => convolution3D_CP_3189_elements(95)); -- 
    cr_3961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(95), ack => RPIPE_maxpool_input_pipe_1387_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1387_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Sample/rr
      -- 
    ca_3962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1387_inst_ack_1, ack => convolution3D_CP_3189_elements(96)); -- 
    rr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(96), ack => type_cast_1391_inst_req_0); -- 
    rr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(96), ack => RPIPE_maxpool_input_pipe_1405_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Sample/ra
      -- 
    ra_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_0, ack => convolution3D_CP_3189_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	319 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Update/ca
      -- 
    ca_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_1, ack => convolution3D_CP_3189_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_update_start_
      -- CP-element group 99: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Update/cr
      -- 
    ra_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1405_inst_ack_0, ack => convolution3D_CP_3189_elements(99)); -- 
    cr_3989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(99), ack => RPIPE_maxpool_input_pipe_1405_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1405_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Sample/rr
      -- 
    ca_3990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1405_inst_ack_1, ack => convolution3D_CP_3189_elements(100)); -- 
    rr_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(100), ack => type_cast_1409_inst_req_0); -- 
    rr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(100), ack => RPIPE_maxpool_input_pipe_1423_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Sample/ra
      -- 
    ra_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1409_inst_ack_0, ack => convolution3D_CP_3189_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	319 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Update/ca
      -- 
    ca_4004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1409_inst_ack_1, ack => convolution3D_CP_3189_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_update_start_
      -- CP-element group 103: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Update/cr
      -- 
    ra_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1423_inst_ack_0, ack => convolution3D_CP_3189_elements(103)); -- 
    cr_4017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(103), ack => RPIPE_maxpool_input_pipe_1423_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	107 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1423_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Sample/rr
      -- 
    ca_4018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1423_inst_ack_1, ack => convolution3D_CP_3189_elements(104)); -- 
    rr_4026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(104), ack => type_cast_1427_inst_req_0); -- 
    rr_4040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(104), ack => RPIPE_maxpool_input_pipe_1441_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Sample/ra
      -- 
    ra_4027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_0, ack => convolution3D_CP_3189_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	319 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Update/ca
      -- 
    ca_4032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_1, ack => convolution3D_CP_3189_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Update/cr
      -- 
    ra_4041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1441_inst_ack_0, ack => convolution3D_CP_3189_elements(107)); -- 
    cr_4045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(107), ack => RPIPE_maxpool_input_pipe_1441_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1441_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Sample/rr
      -- 
    ca_4046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1441_inst_ack_1, ack => convolution3D_CP_3189_elements(108)); -- 
    rr_4054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(108), ack => type_cast_1445_inst_req_0); -- 
    rr_4068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(108), ack => RPIPE_maxpool_input_pipe_1459_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Sample/ra
      -- 
    ra_4055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_0, ack => convolution3D_CP_3189_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	319 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Update/ca
      -- 
    ca_4060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_1, ack => convolution3D_CP_3189_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Update/cr
      -- 
    ra_4069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1459_inst_ack_0, ack => convolution3D_CP_3189_elements(111)); -- 
    cr_4073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(111), ack => RPIPE_maxpool_input_pipe_1459_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1459_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_sample_start_
      -- 
    ca_4074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1459_inst_ack_1, ack => convolution3D_CP_3189_elements(112)); -- 
    rr_4082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(112), ack => type_cast_1463_inst_req_0); -- 
    rr_4096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(112), ack => RPIPE_maxpool_input_pipe_1477_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Sample/$exit
      -- 
    ra_4083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_0, ack => convolution3D_CP_3189_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	319 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_update_completed_
      -- 
    ca_4088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_1, ack => convolution3D_CP_3189_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_update_start_
      -- CP-element group 115: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_sample_completed_
      -- 
    ra_4097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1477_inst_ack_0, ack => convolution3D_CP_3189_elements(115)); -- 
    cr_4101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(115), ack => RPIPE_maxpool_input_pipe_1477_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	119 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1477_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_sample_start_
      -- 
    ca_4102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1477_inst_ack_1, ack => convolution3D_CP_3189_elements(116)); -- 
    rr_4110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(116), ack => type_cast_1481_inst_req_0); -- 
    rr_4124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(116), ack => RPIPE_maxpool_input_pipe_1495_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Sample/$exit
      -- 
    ra_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1481_inst_ack_0, ack => convolution3D_CP_3189_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	319 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Update/ca
      -- 
    ca_4116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1481_inst_ack_1, ack => convolution3D_CP_3189_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_update_start_
      -- CP-element group 119: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_sample_completed_
      -- 
    ra_4125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1495_inst_ack_0, ack => convolution3D_CP_3189_elements(119)); -- 
    cr_4129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(119), ack => RPIPE_maxpool_input_pipe_1495_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1495_update_completed_
      -- 
    ca_4130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1495_inst_ack_1, ack => convolution3D_CP_3189_elements(120)); -- 
    rr_4138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(120), ack => type_cast_1499_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Sample/ra
      -- CP-element group 121: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_sample_completed_
      -- 
    ra_4139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1499_inst_ack_0, ack => convolution3D_CP_3189_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	319 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Update/ca
      -- CP-element group 122: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_update_completed_
      -- 
    ca_4144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1499_inst_ack_1, ack => convolution3D_CP_3189_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	122 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	106 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/ptr_deref_1507_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/ptr_deref_1507_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/ptr_deref_1507_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/word_access_start/word_0/rr
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/ptr_deref_1507_Split/split_ack
      -- 
    rr_4182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(123), ack => ptr_deref_1507_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(110) & convolution3D_CP_3189_elements(122) & convolution3D_CP_3189_elements(114) & convolution3D_CP_3189_elements(118) & convolution3D_CP_3189_elements(90) & convolution3D_CP_3189_elements(94) & convolution3D_CP_3189_elements(98) & convolution3D_CP_3189_elements(102) & convolution3D_CP_3189_elements(106);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/word_access_start/word_0/ra
      -- CP-element group 124: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Sample/word_access_start/$exit
      -- 
    ra_4183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1507_store_0_ack_0, ack => convolution3D_CP_3189_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	319 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/word_access_complete/word_0/ca
      -- CP-element group 125: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/$exit
      -- 
    ca_4194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1507_store_0_ack_1, ack => convolution3D_CP_3189_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: 	87 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520__exit__
      -- CP-element group 126: 	 branch_block_stmt_1049/if_stmt_1521__entry__
      -- CP-element group 126: 	 branch_block_stmt_1049/if_stmt_1521_else_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_1049/R_exitcond28_1522_place
      -- CP-element group 126: 	 branch_block_stmt_1049/if_stmt_1521_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_1049/if_stmt_1521_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_1049/if_stmt_1521_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_1049/if_stmt_1521_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/$exit
      -- CP-element group 126: 	 branch_block_stmt_1049/if_stmt_1521_dead_link/$entry
      -- 
    branch_req_4202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(126), ack => if_stmt_1521_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(125) & convolution3D_CP_3189_elements(87);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	321 
    -- CP-element group 127: 	322 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_1049/assign_stmt_1534_to_assign_stmt_1549__entry__
      -- CP-element group 127: 	 branch_block_stmt_1049/assign_stmt_1534_to_assign_stmt_1549__exit__
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_1049/merge_stmt_1527__exit__
      -- CP-element group 127: 	 branch_block_stmt_1049/assign_stmt_1534_to_assign_stmt_1549/$exit
      -- CP-element group 127: 	 branch_block_stmt_1049/assign_stmt_1534_to_assign_stmt_1549/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/if_stmt_1521_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_1049/if_stmt_1521_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_1049/merge_stmt_1527_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_1049/merge_stmt_1527_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/merge_stmt_1527_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_1049/merge_stmt_1527_PhiAck/dummy
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1521_branch_ack_1, ack => convolution3D_CP_3189_elements(127)); -- 
    rr_5753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(127), ack => type_cast_1555_inst_req_0); -- 
    cr_5758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(127), ack => type_cast_1555_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	315 
    -- CP-element group 128: 	316 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_1049/if_stmt_1521_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_1049/if_stmt_1521_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/$entry
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/$entry
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1521_branch_ack_0, ack => convolution3D_CP_3189_elements(128)); -- 
    rr_5699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(128), ack => type_cast_1364_inst_req_0); -- 
    cr_5704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(128), ack => type_cast_1364_inst_req_1); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	325 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	344 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_1049/if_stmt_1572_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_1049/if_stmt_1572_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_1049/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_1049/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_1049/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_4232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1572_branch_ack_1, ack => convolution3D_CP_3189_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	325 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	326 
    -- CP-element group 130: 	327 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_1049/merge_stmt_1578__exit__
      -- CP-element group 130: 	 branch_block_stmt_1049/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_1049/assign_stmt_1584_to_assign_stmt_1590__entry__
      -- CP-element group 130: 	 branch_block_stmt_1049/assign_stmt_1584_to_assign_stmt_1590__exit__
      -- CP-element group 130: 	 branch_block_stmt_1049/if_stmt_1572_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_1049/if_stmt_1572_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_1049/assign_stmt_1584_to_assign_stmt_1590/$entry
      -- CP-element group 130: 	 branch_block_stmt_1049/assign_stmt_1584_to_assign_stmt_1590/$exit
      -- CP-element group 130: 	 branch_block_stmt_1049/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_1049/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_1049/merge_stmt_1578_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_1049/merge_stmt_1578_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_1049/merge_stmt_1578_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_1049/merge_stmt_1578_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/$entry
      -- CP-element group 130: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/$entry
      -- CP-element group 130: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$entry
      -- 
    else_choice_transition_4236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1572_branch_ack_0, ack => convolution3D_CP_3189_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	339 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_update_start_
      -- 
    ra_4253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1621_inst_ack_0, ack => convolution3D_CP_3189_elements(131)); -- 
    cr_4257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(131), ack => RPIPE_maxpool_input_pipe_1621_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_update_completed_
      -- 
    ca_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1621_inst_ack_1, ack => convolution3D_CP_3189_elements(132)); -- 
    rr_4266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(132), ack => type_cast_1625_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_sample_completed_
      -- 
    ra_4267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_0, ack => convolution3D_CP_3189_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	339 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_update_completed_
      -- 
    ca_4272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_1, ack => convolution3D_CP_3189_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	339 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_sample_completed_
      -- 
    ra_4281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1640_inst_ack_0, ack => convolution3D_CP_3189_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	339 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_update_completed_
      -- 
    ca_4286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1640_inst_ack_1, ack => convolution3D_CP_3189_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646__exit__
      -- CP-element group 137: 	 branch_block_stmt_1049/if_stmt_1647__entry__
      -- CP-element group 137: 	 branch_block_stmt_1049/R_cmpx_xi_1648_place
      -- CP-element group 137: 	 branch_block_stmt_1049/if_stmt_1647_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_1049/if_stmt_1647_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/$exit
      -- CP-element group 137: 	 branch_block_stmt_1049/if_stmt_1647_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1049/if_stmt_1647_else_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1049/if_stmt_1647_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1049/if_stmt_1647_eval_test/branch_req
      -- 
    branch_req_4294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(137), ack => if_stmt_1647_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(134) & convolution3D_CP_3189_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	329 
    -- CP-element group 138: 	330 
    -- CP-element group 138: 	332 
    -- CP-element group 138: 	333 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_1049/if_stmt_1647_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_1049/if_stmt_1647_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1647_branch_ack_1, ack => convolution3D_CP_3189_elements(138)); -- 
    rr_5815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(138), ack => type_cast_1599_inst_req_0); -- 
    cr_5820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(138), ack => type_cast_1599_inst_req_1); -- 
    rr_5838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(138), ack => type_cast_1606_inst_req_0); -- 
    cr_5843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(138), ack => type_cast_1606_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	340 
    -- CP-element group 139: 	341 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_1049/if_stmt_1647_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_1049/if_stmt_1647_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/$entry
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/$entry
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1647_branch_ack_0, ack => convolution3D_CP_3189_elements(139)); -- 
    rr_5874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(139), ack => type_cast_1657_inst_req_0); -- 
    cr_5879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(139), ack => type_cast_1657_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	343 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_sample_complete
      -- CP-element group 140: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Sample/$exit
      -- 
    ack_4334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1686_index_offset_ack_0, ack => convolution3D_CP_3189_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	343 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_request/req
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Update/$exit
      -- 
    ack_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1686_index_offset_ack_1, ack => convolution3D_CP_3189_elements(141)); -- 
    req_4348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(141), ack => addr_of_1687_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_request/ack
      -- CP-element group 142: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_request/$exit
      -- 
    ack_4349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1687_final_reg_ack_0, ack => convolution3D_CP_3189_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	343 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/word_access_start/word_0/rr
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/ptr_deref_1690_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/ptr_deref_1690_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/ptr_deref_1690_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/ptr_deref_1690_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_word_addrgen/root_register_ack
      -- 
    ack_4354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1687_final_reg_ack_1, ack => convolution3D_CP_3189_elements(143)); -- 
    rr_4392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(143), ack => ptr_deref_1690_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/word_access_start/word_0/ra
      -- CP-element group 144: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Sample/$exit
      -- 
    ra_4393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1690_store_0_ack_0, ack => convolution3D_CP_3189_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	343 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/word_access_complete/word_0/ca
      -- CP-element group 145: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/word_access_complete/word_0/$exit
      -- 
    ca_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1690_store_0_ack_1, ack => convolution3D_CP_3189_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	140 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	344 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692__exit__
      -- CP-element group 146: 	 branch_block_stmt_1049/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/$exit
      -- CP-element group 146: 	 branch_block_stmt_1049/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_1049/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(140) & convolution3D_CP_3189_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	344 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_sample_completed_
      -- 
    ra_4416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1697_inst_ack_0, ack => convolution3D_CP_3189_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	344 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_update_completed_
      -- 
    ca_4421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1697_inst_ack_1, ack => convolution3D_CP_3189_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	344 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Sample/$exit
      -- 
    ra_4430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_0, ack => convolution3D_CP_3189_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	344 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Update/$exit
      -- 
    ca_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_1, ack => convolution3D_CP_3189_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	344 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Sample/$exit
      -- 
    ra_4444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1705_inst_ack_0, ack => convolution3D_CP_3189_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	344 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Update/$exit
      -- 
    ca_4449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1705_inst_ack_1, ack => convolution3D_CP_3189_elements(152)); -- 
    -- CP-element group 153:  branch  join  transition  place  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: 	152 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (10) 
      -- CP-element group 153: 	 branch_block_stmt_1049/R_cmp161379_1744_place
      -- CP-element group 153: 	 branch_block_stmt_1049/if_stmt_1743__entry__
      -- CP-element group 153: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742__exit__
      -- CP-element group 153: 	 branch_block_stmt_1049/if_stmt_1743_dead_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_1049/if_stmt_1743_else_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_1049/if_stmt_1743_if_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/$exit
      -- CP-element group 153: 	 branch_block_stmt_1049/if_stmt_1743_eval_test/branch_req
      -- CP-element group 153: 	 branch_block_stmt_1049/if_stmt_1743_eval_test/$entry
      -- CP-element group 153: 	 branch_block_stmt_1049/if_stmt_1743_eval_test/$exit
      -- 
    branch_req_4457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(153), ack => if_stmt_1743_branch_req_0); -- 
    convolution3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(150) & convolution3D_CP_3189_elements(152) & convolution3D_CP_3189_elements(148);
      gj_convolution3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	159 
    -- CP-element group 154: 	160 
    -- CP-element group 154: 	161 
    -- CP-element group 154: 	164 
    -- CP-element group 154: 	156 
    -- CP-element group 154: 	157 
    -- CP-element group 154: 	158 
    -- CP-element group 154: 	166 
    -- CP-element group 154:  members (36) 
      -- CP-element group 154: 	 branch_block_stmt_1049/merge_stmt_1749__exit__
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816__entry__
      -- CP-element group 154: 	 branch_block_stmt_1049/ifx_xend_bbx_xnph
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1049/if_stmt_1743_if_link/if_choice_transition
      -- CP-element group 154: 	 branch_block_stmt_1049/if_stmt_1743_if_link/$exit
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1049/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 154: 	 branch_block_stmt_1049/merge_stmt_1749_PhiReqMerge
      -- CP-element group 154: 	 branch_block_stmt_1049/merge_stmt_1749_PhiAck/$entry
      -- CP-element group 154: 	 branch_block_stmt_1049/merge_stmt_1749_PhiAck/$exit
      -- CP-element group 154: 	 branch_block_stmt_1049/merge_stmt_1749_PhiAck/dummy
      -- 
    if_choice_transition_4462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1743_branch_ack_1, ack => convolution3D_CP_3189_elements(154)); -- 
    rr_4507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1782_inst_req_0); -- 
    cr_4512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1782_inst_req_1); -- 
    rr_4493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1773_inst_req_0); -- 
    cr_4484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1764_inst_req_1); -- 
    cr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1773_inst_req_1); -- 
    rr_4479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1764_inst_req_0); -- 
    cr_4526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1791_inst_req_1); -- 
    cr_4540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(154), ack => type_cast_1796_inst_req_1); -- 
    -- CP-element group 155:  transition  place  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	354 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1049/ifx_xend_forx_xend215
      -- CP-element group 155: 	 branch_block_stmt_1049/if_stmt_1743_else_link/else_choice_transition
      -- CP-element group 155: 	 branch_block_stmt_1049/if_stmt_1743_else_link/$exit
      -- CP-element group 155: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/$entry
      -- CP-element group 155: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/phi_stmt_2013/$entry
      -- CP-element group 155: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/$entry
      -- 
    else_choice_transition_4466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1743_branch_ack_0, ack => convolution3D_CP_3189_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_sample_completed_
      -- 
    ra_4480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_0, ack => convolution3D_CP_3189_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1764_update_completed_
      -- 
    ca_4485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_1, ack => convolution3D_CP_3189_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Sample/ra
      -- 
    ra_4494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_0, ack => convolution3D_CP_3189_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	154 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1773_Update/ca
      -- 
    ca_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_1, ack => convolution3D_CP_3189_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	154 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Sample/ra
      -- 
    ra_4508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1782_inst_ack_0, ack => convolution3D_CP_3189_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	154 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1782_Update/ca
      -- 
    ca_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1782_inst_ack_1, ack => convolution3D_CP_3189_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	159 
    -- CP-element group 162: 	161 
    -- CP-element group 162: 	157 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Sample/rr
      -- 
    rr_4521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(162), ack => type_cast_1791_inst_req_0); -- 
    convolution3D_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(159) & convolution3D_CP_3189_elements(161) & convolution3D_CP_3189_elements(157);
      gj_convolution3D_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Sample/ra
      -- 
    ra_4522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_0, ack => convolution3D_CP_3189_elements(163)); -- 
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	154 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1791_Update/ca
      -- CP-element group 164: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Sample/rr
      -- 
    ca_4527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_1, ack => convolution3D_CP_3189_elements(164)); -- 
    rr_4535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(164), ack => type_cast_1796_inst_req_0); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Sample/ra
      -- 
    ra_4536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1796_inst_ack_0, ack => convolution3D_CP_3189_elements(165)); -- 
    -- CP-element group 166:  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	154 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	345 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816__exit__
      -- CP-element group 166: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163
      -- CP-element group 166: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/$exit
      -- CP-element group 166: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_1049/assign_stmt_1755_to_assign_stmt_1816/type_cast_1796_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1819/$entry
      -- CP-element group 166: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$entry
      -- 
    ca_4541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1796_inst_ack_1, ack => convolution3D_CP_3189_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	350 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	206 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_sample_complete
      -- CP-element group 167: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Sample/ack
      -- 
    ack_4570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1831_index_offset_ack_0, ack => convolution3D_CP_3189_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	350 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (11) 
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_offset_calculated
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Update/ack
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_base_plus_offset/$entry
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_base_plus_offset/$exit
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_request/$entry
      -- CP-element group 168: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_request/req
      -- 
    ack_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1831_index_offset_ack_1, ack => convolution3D_CP_3189_elements(168)); -- 
    req_4584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(168), ack => addr_of_1832_final_reg_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_request/$exit
      -- CP-element group 169: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_request/ack
      -- 
    ack_4585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1832_final_reg_ack_0, ack => convolution3D_CP_3189_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	350 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	203 
    -- CP-element group 170:  members (19) 
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_complete/$exit
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_complete/ack
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_word_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_address_resized
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_addr_resize/$entry
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_addr_resize/$exit
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_addr_resize/base_resize_req
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_addr_resize/base_resize_ack
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_word_addrgen/$entry
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_word_addrgen/$exit
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_word_addrgen/root_register_req
      -- CP-element group 170: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_word_addrgen/root_register_ack
      -- 
    ack_4590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1832_final_reg_ack_1, ack => convolution3D_CP_3189_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	350 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_update_start_
      -- CP-element group 171: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Sample/ra
      -- CP-element group 171: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Update/cr
      -- 
    ra_4599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1835_inst_ack_0, ack => convolution3D_CP_3189_elements(171)); -- 
    cr_4603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(171), ack => RPIPE_maxpool_input_pipe_1835_inst_req_1); -- 
    -- CP-element group 172:  fork  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: 	175 
    -- CP-element group 172:  members (9) 
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Sample/rr
      -- 
    ca_4604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1835_inst_ack_1, ack => convolution3D_CP_3189_elements(172)); -- 
    rr_4612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(172), ack => type_cast_1839_inst_req_0); -- 
    rr_4626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(172), ack => RPIPE_maxpool_input_pipe_1848_inst_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Sample/ra
      -- 
    ra_4613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1839_inst_ack_0, ack => convolution3D_CP_3189_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	350 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	203 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Update/ca
      -- 
    ca_4618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1839_inst_ack_1, ack => convolution3D_CP_3189_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	172 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Update/cr
      -- 
    ra_4627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1848_inst_ack_0, ack => convolution3D_CP_3189_elements(175)); -- 
    cr_4631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(175), ack => RPIPE_maxpool_input_pipe_1848_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1848_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Sample/rr
      -- 
    ca_4632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1848_inst_ack_1, ack => convolution3D_CP_3189_elements(176)); -- 
    rr_4640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(176), ack => type_cast_1852_inst_req_0); -- 
    rr_4654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(176), ack => RPIPE_maxpool_input_pipe_1866_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Sample/ra
      -- 
    ra_4641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1852_inst_ack_0, ack => convolution3D_CP_3189_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	350 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	203 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Update/ca
      -- 
    ca_4646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1852_inst_ack_1, ack => convolution3D_CP_3189_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Update/cr
      -- 
    ra_4655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1866_inst_ack_0, ack => convolution3D_CP_3189_elements(179)); -- 
    cr_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(179), ack => RPIPE_maxpool_input_pipe_1866_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1866_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Sample/rr
      -- 
    ca_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1866_inst_ack_1, ack => convolution3D_CP_3189_elements(180)); -- 
    rr_4668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(180), ack => type_cast_1870_inst_req_0); -- 
    rr_4682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(180), ack => RPIPE_maxpool_input_pipe_1884_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Sample/ra
      -- 
    ra_4669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1870_inst_ack_0, ack => convolution3D_CP_3189_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	350 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	203 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Update/ca
      -- 
    ca_4674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1870_inst_ack_1, ack => convolution3D_CP_3189_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_update_start_
      -- CP-element group 183: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Update/cr
      -- 
    ra_4683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1884_inst_ack_0, ack => convolution3D_CP_3189_elements(183)); -- 
    cr_4687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(183), ack => RPIPE_maxpool_input_pipe_1884_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1884_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Sample/rr
      -- 
    ca_4688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1884_inst_ack_1, ack => convolution3D_CP_3189_elements(184)); -- 
    rr_4696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(184), ack => type_cast_1888_inst_req_0); -- 
    rr_4710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(184), ack => RPIPE_maxpool_input_pipe_1902_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Sample/ra
      -- 
    ra_4697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_0, ack => convolution3D_CP_3189_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	350 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	203 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Update/ca
      -- 
    ca_4702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_1, ack => convolution3D_CP_3189_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_update_start_
      -- CP-element group 187: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Update/cr
      -- 
    ra_4711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1902_inst_ack_0, ack => convolution3D_CP_3189_elements(187)); -- 
    cr_4715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(187), ack => RPIPE_maxpool_input_pipe_1902_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1902_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Sample/rr
      -- 
    ca_4716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1902_inst_ack_1, ack => convolution3D_CP_3189_elements(188)); -- 
    rr_4724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(188), ack => type_cast_1906_inst_req_0); -- 
    rr_4738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(188), ack => RPIPE_maxpool_input_pipe_1920_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Sample/ra
      -- 
    ra_4725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1906_inst_ack_0, ack => convolution3D_CP_3189_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	350 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	203 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Update/ca
      -- 
    ca_4730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1906_inst_ack_1, ack => convolution3D_CP_3189_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_update_start_
      -- CP-element group 191: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Update/cr
      -- 
    ra_4739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1920_inst_ack_0, ack => convolution3D_CP_3189_elements(191)); -- 
    cr_4743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(191), ack => RPIPE_maxpool_input_pipe_1920_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1920_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Sample/rr
      -- 
    ca_4744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1920_inst_ack_1, ack => convolution3D_CP_3189_elements(192)); -- 
    rr_4752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(192), ack => type_cast_1924_inst_req_0); -- 
    rr_4766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(192), ack => RPIPE_maxpool_input_pipe_1938_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Sample/ra
      -- 
    ra_4753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1924_inst_ack_0, ack => convolution3D_CP_3189_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	350 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	203 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Update/ca
      -- 
    ca_4758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1924_inst_ack_1, ack => convolution3D_CP_3189_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_update_start_
      -- CP-element group 195: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Update/cr
      -- 
    ra_4767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1938_inst_ack_0, ack => convolution3D_CP_3189_elements(195)); -- 
    cr_4771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(195), ack => RPIPE_maxpool_input_pipe_1938_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1938_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Sample/rr
      -- 
    ca_4772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1938_inst_ack_1, ack => convolution3D_CP_3189_elements(196)); -- 
    rr_4780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(196), ack => type_cast_1942_inst_req_0); -- 
    rr_4794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(196), ack => RPIPE_maxpool_input_pipe_1956_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Sample/ra
      -- 
    ra_4781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1942_inst_ack_0, ack => convolution3D_CP_3189_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	350 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	203 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Update/ca
      -- 
    ca_4786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1942_inst_ack_1, ack => convolution3D_CP_3189_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_update_start_
      -- CP-element group 199: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Update/cr
      -- 
    ra_4795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1956_inst_ack_0, ack => convolution3D_CP_3189_elements(199)); -- 
    cr_4799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(199), ack => RPIPE_maxpool_input_pipe_1956_inst_req_1); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1956_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Sample/rr
      -- 
    ca_4800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1956_inst_ack_1, ack => convolution3D_CP_3189_elements(200)); -- 
    rr_4808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(200), ack => type_cast_1960_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Sample/ra
      -- 
    ra_4809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1960_inst_ack_0, ack => convolution3D_CP_3189_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	350 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Update/ca
      -- 
    ca_4814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1960_inst_ack_1, ack => convolution3D_CP_3189_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	174 
    -- CP-element group 203: 	178 
    -- CP-element group 203: 	186 
    -- CP-element group 203: 	170 
    -- CP-element group 203: 	190 
    -- CP-element group 203: 	198 
    -- CP-element group 203: 	182 
    -- CP-element group 203: 	194 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/ptr_deref_1968_Split/$entry
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/ptr_deref_1968_Split/$exit
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/ptr_deref_1968_Split/split_req
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/ptr_deref_1968_Split/split_ack
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/word_access_start/$entry
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/word_access_start/word_0/$entry
      -- CP-element group 203: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/word_access_start/word_0/rr
      -- 
    rr_4852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(203), ack => ptr_deref_1968_store_0_req_0); -- 
    convolution3D_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(174) & convolution3D_CP_3189_elements(178) & convolution3D_CP_3189_elements(186) & convolution3D_CP_3189_elements(170) & convolution3D_CP_3189_elements(190) & convolution3D_CP_3189_elements(198) & convolution3D_CP_3189_elements(182) & convolution3D_CP_3189_elements(194) & convolution3D_CP_3189_elements(202);
      gj_convolution3D_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/word_access_start/$exit
      -- CP-element group 204: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/word_access_start/word_0/$exit
      -- CP-element group 204: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Sample/word_access_start/word_0/ra
      -- 
    ra_4853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_store_0_ack_0, ack => convolution3D_CP_3189_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	350 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/word_access_complete/$exit
      -- CP-element group 205: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/word_access_complete/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/word_access_complete/word_0/ca
      -- 
    ca_4864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_store_0_ack_1, ack => convolution3D_CP_3189_elements(205)); -- 
    -- CP-element group 206:  branch  join  transition  place  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	167 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (10) 
      -- CP-element group 206: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981__exit__
      -- CP-element group 206: 	 branch_block_stmt_1049/if_stmt_1982__entry__
      -- CP-element group 206: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/$exit
      -- CP-element group 206: 	 branch_block_stmt_1049/if_stmt_1982_dead_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_1049/if_stmt_1982_eval_test/$entry
      -- CP-element group 206: 	 branch_block_stmt_1049/if_stmt_1982_eval_test/$exit
      -- CP-element group 206: 	 branch_block_stmt_1049/if_stmt_1982_eval_test/branch_req
      -- CP-element group 206: 	 branch_block_stmt_1049/R_exitcond_1983_place
      -- CP-element group 206: 	 branch_block_stmt_1049/if_stmt_1982_if_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_1049/if_stmt_1982_else_link/$entry
      -- 
    branch_req_4872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(206), ack => if_stmt_1982_branch_req_0); -- 
    convolution3D_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(167) & convolution3D_CP_3189_elements(205);
      gj_convolution3D_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	351 
    -- CP-element group 207: 	352 
    -- CP-element group 207:  members (24) 
      -- CP-element group 207: 	 branch_block_stmt_1049/merge_stmt_1988__exit__
      -- CP-element group 207: 	 branch_block_stmt_1049/assign_stmt_1995_to_assign_stmt_2010__entry__
      -- CP-element group 207: 	 branch_block_stmt_1049/assign_stmt_1995_to_assign_stmt_2010__exit__
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 207: 	 branch_block_stmt_1049/if_stmt_1982_if_link/$exit
      -- CP-element group 207: 	 branch_block_stmt_1049/if_stmt_1982_if_link/if_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 207: 	 branch_block_stmt_1049/assign_stmt_1995_to_assign_stmt_2010/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/assign_stmt_1995_to_assign_stmt_2010/$exit
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_1049/merge_stmt_1988_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_1049/merge_stmt_1988_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/merge_stmt_1988_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_1049/merge_stmt_1988_PhiAck/dummy
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1982_branch_ack_1, ack => convolution3D_CP_3189_elements(207)); -- 
    rr_5982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(207), ack => type_cast_2016_inst_req_0); -- 
    cr_5987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(207), ack => type_cast_2016_inst_req_1); -- 
    -- CP-element group 208:  fork  transition  place  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	346 
    -- CP-element group 208: 	347 
    -- CP-element group 208:  members (12) 
      -- CP-element group 208: 	 branch_block_stmt_1049/if_stmt_1982_else_link/$exit
      -- CP-element group 208: 	 branch_block_stmt_1049/if_stmt_1982_else_link/else_choice_transition
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/$entry
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$entry
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/$entry
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/$entry
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1982_branch_ack_0, ack => convolution3D_CP_3189_elements(208)); -- 
    rr_5939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(208), ack => type_cast_1822_inst_req_0); -- 
    cr_5944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(208), ack => type_cast_1822_inst_req_1); -- 
    -- CP-element group 209:  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	356 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	375 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_1049/if_stmt_2033_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_1049/if_stmt_2033_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_1049/forx_xend215_ifx_xend227
      -- CP-element group 209: 	 branch_block_stmt_1049/forx_xend215_ifx_xend227_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_1049/forx_xend215_ifx_xend227_PhiReq/$exit
      -- 
    if_choice_transition_4902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2033_branch_ack_1, ack => convolution3D_CP_3189_elements(209)); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	356 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (18) 
      -- CP-element group 210: 	 branch_block_stmt_1049/merge_stmt_2039__exit__
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055__entry__
      -- CP-element group 210: 	 branch_block_stmt_1049/if_stmt_2033_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_1049/if_stmt_2033_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_1049/forx_xend215_bbx_xnphx_xi356
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/$entry
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_update_start_
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_1049/forx_xend215_bbx_xnphx_xi356_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_1049/forx_xend215_bbx_xnphx_xi356_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_1049/merge_stmt_2039_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_1049/merge_stmt_2039_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_1049/merge_stmt_2039_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_1049/merge_stmt_2039_PhiAck/dummy
      -- 
    else_choice_transition_4906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2033_branch_ack_0, ack => convolution3D_CP_3189_elements(210)); -- 
    rr_4919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(210), ack => type_cast_2048_inst_req_0); -- 
    cr_4924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(210), ack => type_cast_2048_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Sample/ra
      -- 
    ra_4920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_0, ack => convolution3D_CP_3189_elements(211)); -- 
    -- CP-element group 212:  fork  transition  place  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	357 
    -- CP-element group 212: 	358 
    -- CP-element group 212:  members (11) 
      -- CP-element group 212: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055__exit__
      -- CP-element group 212: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365
      -- CP-element group 212: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/$exit
      -- CP-element group 212: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_1049/assign_stmt_2045_to_assign_stmt_2055/type_cast_2048_Update/ca
      -- CP-element group 212: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/$entry
      -- CP-element group 212: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/$entry
      -- CP-element group 212: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$entry
      -- 
    ca_4925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_1, ack => convolution3D_CP_3189_elements(212)); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	370 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_update_start_
      -- CP-element group 213: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Sample/ra
      -- CP-element group 213: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Update/cr
      -- 
    ra_4937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2086_inst_ack_0, ack => convolution3D_CP_3189_elements(213)); -- 
    cr_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(213), ack => RPIPE_maxpool_input_pipe_2086_inst_req_1); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Update/ca
      -- CP-element group 214: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Sample/rr
      -- 
    ca_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2086_inst_ack_1, ack => convolution3D_CP_3189_elements(214)); -- 
    rr_4950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(214), ack => type_cast_2090_inst_req_0); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Sample/ra
      -- 
    ra_4951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2090_inst_ack_0, ack => convolution3D_CP_3189_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	370 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	219 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Update/ca
      -- 
    ca_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2090_inst_ack_1, ack => convolution3D_CP_3189_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	370 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Sample/ra
      -- 
    ra_4965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2105_inst_ack_0, ack => convolution3D_CP_3189_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	370 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Update/ca
      -- 
    ca_4970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2105_inst_ack_1, ack => convolution3D_CP_3189_elements(218)); -- 
    -- CP-element group 219:  branch  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	216 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (10) 
      -- CP-element group 219: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111__exit__
      -- CP-element group 219: 	 branch_block_stmt_1049/if_stmt_2112__entry__
      -- CP-element group 219: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/$exit
      -- CP-element group 219: 	 branch_block_stmt_1049/if_stmt_2112_dead_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_1049/if_stmt_2112_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_1049/if_stmt_2112_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_1049/if_stmt_2112_eval_test/branch_req
      -- CP-element group 219: 	 branch_block_stmt_1049/R_cmpx_xi364_2113_place
      -- CP-element group 219: 	 branch_block_stmt_1049/if_stmt_2112_if_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_1049/if_stmt_2112_else_link/$entry
      -- 
    branch_req_4978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(219), ack => if_stmt_2112_branch_req_0); -- 
    convolution3D_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(216) & convolution3D_CP_3189_elements(218);
      gj_convolution3D_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  place  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	360 
    -- CP-element group 220: 	361 
    -- CP-element group 220: 	363 
    -- CP-element group 220: 	364 
    -- CP-element group 220:  members (20) 
      -- CP-element group 220: 	 branch_block_stmt_1049/if_stmt_2112_if_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_1049/if_stmt_2112_if_link/if_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Update/cr
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2112_branch_ack_1, ack => convolution3D_CP_3189_elements(220)); -- 
    rr_6055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(220), ack => type_cast_2068_inst_req_0); -- 
    cr_6060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(220), ack => type_cast_2068_inst_req_1); -- 
    rr_6078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(220), ack => type_cast_2061_inst_req_0); -- 
    cr_6083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(220), ack => type_cast_2061_inst_req_1); -- 
    -- CP-element group 221:  fork  transition  place  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	371 
    -- CP-element group 221: 	372 
    -- CP-element group 221:  members (12) 
      -- CP-element group 221: 	 branch_block_stmt_1049/if_stmt_2112_else_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_1049/if_stmt_2112_else_link/else_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/$entry
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/$entry
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/$entry
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Sample/rr
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2112_branch_ack_0, ack => convolution3D_CP_3189_elements(221)); -- 
    rr_6114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(221), ack => type_cast_2122_inst_req_0); -- 
    cr_6119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(221), ack => type_cast_2122_inst_req_1); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	374 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Sample/ack
      -- 
    ack_5018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2151_index_offset_ack_0, ack => convolution3D_CP_3189_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	374 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_request/req
      -- 
    ack_5023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2151_index_offset_ack_1, ack => convolution3D_CP_3189_elements(223)); -- 
    req_5032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(223), ack => addr_of_2152_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_request/ack
      -- 
    ack_5033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2152_final_reg_ack_0, ack => convolution3D_CP_3189_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	374 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/ptr_deref_2155_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/ptr_deref_2155_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/ptr_deref_2155_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/ptr_deref_2155_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/word_access_start/word_0/rr
      -- 
    ack_5038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2152_final_reg_ack_1, ack => convolution3D_CP_3189_elements(225)); -- 
    rr_5076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(225), ack => ptr_deref_2155_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Sample/word_access_start/word_0/ra
      -- 
    ra_5077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2155_store_0_ack_0, ack => convolution3D_CP_3189_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	374 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/word_access_complete/word_0/ca
      -- 
    ca_5088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2155_store_0_ack_1, ack => convolution3D_CP_3189_elements(227)); -- 
    -- CP-element group 228:  join  transition  place  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: 	222 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	375 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157__exit__
      -- CP-element group 228: 	 branch_block_stmt_1049/getRemainingElementsx_xexit373_ifx_xend227
      -- CP-element group 228: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/$exit
      -- CP-element group 228: 	 branch_block_stmt_1049/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_1049/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(227) & convolution3D_CP_3189_elements(222);
      gj_convolution3D_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	376 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (5) 
      -- CP-element group 229: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_sample_completed_
      -- CP-element group 229: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/word_access_start/$exit
      -- CP-element group 229: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/word_access_start/word_0/$exit
      -- CP-element group 229: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/word_access_start/word_0/ra
      -- 
    ra_5130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2169_store_0_ack_0, ack => convolution3D_CP_3189_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	376 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230: 	232 
    -- CP-element group 230: 	233 
    -- CP-element group 230:  members (18) 
      -- CP-element group 230: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172__exit__
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184__entry__
      -- CP-element group 230: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/$exit
      -- CP-element group 230: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/word_access_complete/$exit
      -- CP-element group 230: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/word_access_complete/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/word_access_complete/word_0/ca
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/$entry
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_update_start_
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Sample/crr
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Update/ccr
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Sample/req
      -- 
    ca_5141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2169_store_0_ack_1, ack => convolution3D_CP_3189_elements(230)); -- 
    crr_5152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(230), ack => call_stmt_2175_call_req_0); -- 
    ccr_5157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(230), ack => call_stmt_2175_call_req_1); -- 
    req_5166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(230), ack => WPIPE_output_pipe_2176_inst_req_0); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Sample/cra
      -- 
    cra_5153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2175_call_ack_0, ack => convolution3D_CP_3189_elements(231)); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	239 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/call_stmt_2175_Update/cca
      -- 
    cca_5158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2175_call_ack_1, ack => convolution3D_CP_3189_elements(232)); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	230 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_update_start_
      -- CP-element group 233: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Sample/ack
      -- CP-element group 233: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Update/req
      -- 
    ack_5167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2176_inst_ack_0, ack => convolution3D_CP_3189_elements(233)); -- 
    req_5171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(233), ack => WPIPE_output_pipe_2176_inst_req_1); -- 
    -- CP-element group 234:  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2176_Update/ack
      -- CP-element group 234: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Sample/req
      -- 
    ack_5172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2176_inst_ack_1, ack => convolution3D_CP_3189_elements(234)); -- 
    req_5180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(234), ack => WPIPE_output_pipe_2179_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_update_start_
      -- CP-element group 235: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Update/req
      -- 
    ack_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2179_inst_ack_0, ack => convolution3D_CP_3189_elements(235)); -- 
    req_5185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(235), ack => WPIPE_output_pipe_2179_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2179_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Sample/req
      -- 
    ack_5186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2179_inst_ack_1, ack => convolution3D_CP_3189_elements(236)); -- 
    req_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(236), ack => WPIPE_output_pipe_2182_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_update_start_
      -- CP-element group 237: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Update/req
      -- 
    ack_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2182_inst_ack_0, ack => convolution3D_CP_3189_elements(237)); -- 
    req_5199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(237), ack => WPIPE_output_pipe_2182_inst_req_1); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/WPIPE_output_pipe_2182_Update/ack
      -- 
    ack_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2182_inst_ack_1, ack => convolution3D_CP_3189_elements(238)); -- 
    -- CP-element group 239:  join  fork  transition  place  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: 	232 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239: 	241 
    -- CP-element group 239: 	242 
    -- CP-element group 239: 	243 
    -- CP-element group 239:  members (16) 
      -- CP-element group 239: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184__exit__
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215__entry__
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Sample/rr
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_update_start_
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Update/cr
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Update/cr
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_1049/call_stmt_2175_to_assign_stmt_2184/$exit
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/$entry
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_update_start_
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Sample/rr
      -- 
    rr_5225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(239), ack => type_cast_2209_inst_req_0); -- 
    cr_5216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(239), ack => type_cast_2199_inst_req_1); -- 
    cr_5230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(239), ack => type_cast_2209_inst_req_1); -- 
    rr_5211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(239), ack => type_cast_2199_inst_req_0); -- 
    convolution3D_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(238) & convolution3D_CP_3189_elements(232);
      gj_convolution3D_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Sample/ra
      -- 
    ra_5212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => convolution3D_CP_3189_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	244 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Update/ca
      -- CP-element group 241: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2199_update_completed_
      -- 
    ca_5217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_1, ack => convolution3D_CP_3189_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	239 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Sample/ra
      -- CP-element group 242: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_sample_completed_
      -- 
    ra_5226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2209_inst_ack_0, ack => convolution3D_CP_3189_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	239 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Update/ca
      -- CP-element group 243: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/type_cast_2209_Update/$exit
      -- 
    ca_5231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2209_inst_ack_1, ack => convolution3D_CP_3189_elements(243)); -- 
    -- CP-element group 244:  join  transition  place  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	241 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	377 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215__exit__
      -- CP-element group 244: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody
      -- CP-element group 244: 	 branch_block_stmt_1049/assign_stmt_2191_to_assign_stmt_2215/$exit
      -- CP-element group 244: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- CP-element group 244: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2218/$entry
      -- CP-element group 244: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/$entry
      -- 
    convolution3D_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(241) & convolution3D_CP_3189_elements(243);
      gj_convolution3D_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	382 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Update/req
      -- CP-element group 245: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_update_start_
      -- CP-element group 245: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_sample_completed_
      -- 
    ack_5243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2231_inst_ack_0, ack => convolution3D_CP_3189_elements(245)); -- 
    req_5247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(245), ack => WPIPE_num_out_pipe_2231_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_update_completed_
      -- 
    ack_5248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2231_inst_ack_1, ack => convolution3D_CP_3189_elements(246)); -- 
    req_5256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(246), ack => WPIPE_num_out_pipe_2234_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Update/req
      -- CP-element group 247: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_sample_completed_
      -- 
    ack_5257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2234_inst_ack_0, ack => convolution3D_CP_3189_elements(247)); -- 
    req_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(247), ack => WPIPE_num_out_pipe_2234_inst_req_1); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	253 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2234_update_completed_
      -- 
    ack_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2234_inst_ack_1, ack => convolution3D_CP_3189_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	382 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Sample/cra
      -- CP-element group 249: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Sample/$exit
      -- 
    cra_5271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2245_call_ack_0, ack => convolution3D_CP_3189_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	382 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	253 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Update/cca
      -- CP-element group 250: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_update_completed_
      -- 
    cca_5276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2245_call_ack_1, ack => convolution3D_CP_3189_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	382 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Sample/cra
      -- CP-element group 251: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_sample_completed_
      -- 
    cra_5285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2249_call_ack_0, ack => convolution3D_CP_3189_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	382 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Update/cca
      -- CP-element group 252: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_update_completed_
      -- 
    cca_5290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2249_call_ack_1, ack => convolution3D_CP_3189_elements(252)); -- 
    -- CP-element group 253:  branch  join  transition  place  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	248 
    -- CP-element group 253: 	250 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (10) 
      -- CP-element group 253: 	 branch_block_stmt_1049/if_stmt_2261__entry__
      -- CP-element group 253: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260__exit__
      -- CP-element group 253: 	 branch_block_stmt_1049/R_exitcond5_2262_place
      -- CP-element group 253: 	 branch_block_stmt_1049/if_stmt_2261_else_link/$entry
      -- CP-element group 253: 	 branch_block_stmt_1049/if_stmt_2261_if_link/$entry
      -- CP-element group 253: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/$exit
      -- CP-element group 253: 	 branch_block_stmt_1049/if_stmt_2261_eval_test/branch_req
      -- CP-element group 253: 	 branch_block_stmt_1049/if_stmt_2261_eval_test/$exit
      -- CP-element group 253: 	 branch_block_stmt_1049/if_stmt_2261_eval_test/$entry
      -- CP-element group 253: 	 branch_block_stmt_1049/if_stmt_2261_dead_link/$entry
      -- 
    branch_req_5298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(253), ack => if_stmt_2261_branch_req_0); -- 
    convolution3D_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(248) & convolution3D_CP_3189_elements(250) & convolution3D_CP_3189_elements(252);
      gj_convolution3D_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	257 
    -- CP-element group 254: 	258 
    -- CP-element group 254:  members (21) 
      -- CP-element group 254: 	 branch_block_stmt_1049/merge_stmt_2267__exit__
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275__entry__
      -- CP-element group 254: 	 branch_block_stmt_1049/whilex_xbody_whilex_xend
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Sample/rr
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Update/cr
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Sample/rr
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_update_start_
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/$entry
      -- CP-element group 254: 	 branch_block_stmt_1049/if_stmt_2261_if_link/if_choice_transition
      -- CP-element group 254: 	 branch_block_stmt_1049/if_stmt_2261_if_link/$exit
      -- CP-element group 254: 	 branch_block_stmt_1049/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 254: 	 branch_block_stmt_1049/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 254: 	 branch_block_stmt_1049/merge_stmt_2267_PhiReqMerge
      -- CP-element group 254: 	 branch_block_stmt_1049/merge_stmt_2267_PhiAck/$entry
      -- CP-element group 254: 	 branch_block_stmt_1049/merge_stmt_2267_PhiAck/$exit
      -- CP-element group 254: 	 branch_block_stmt_1049/merge_stmt_2267_PhiAck/dummy
      -- 
    if_choice_transition_5303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2261_branch_ack_1, ack => convolution3D_CP_3189_elements(254)); -- 
    rr_5334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(254), ack => RPIPE_input_done_pipe_2274_inst_req_0); -- 
    cr_5325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(254), ack => type_cast_2271_inst_req_1); -- 
    rr_5320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(254), ack => type_cast_2271_inst_req_0); -- 
    -- CP-element group 255:  fork  transition  place  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	378 
    -- CP-element group 255: 	379 
    -- CP-element group 255:  members (12) 
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody
      -- CP-element group 255: 	 branch_block_stmt_1049/if_stmt_2261_else_link/else_choice_transition
      -- CP-element group 255: 	 branch_block_stmt_1049/if_stmt_2261_else_link/$exit
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/$entry
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/$entry
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/$entry
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/$entry
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Sample/rr
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2261_branch_ack_0, ack => convolution3D_CP_3189_elements(255)); -- 
    rr_6167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(255), ack => type_cast_2224_inst_req_0); -- 
    cr_6172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(255), ack => type_cast_2224_inst_req_1); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Sample/ra
      -- CP-element group 256: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_sample_completed_
      -- 
    ra_5321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2271_inst_ack_0, ack => convolution3D_CP_3189_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	254 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	260 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Update/ca
      -- CP-element group 257: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/type_cast_2271_update_completed_
      -- 
    ca_5326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2271_inst_ack_1, ack => convolution3D_CP_3189_elements(257)); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	254 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Update/cr
      -- CP-element group 258: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Sample/ra
      -- CP-element group 258: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_update_start_
      -- CP-element group 258: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_sample_completed_
      -- 
    ra_5335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2274_inst_ack_0, ack => convolution3D_CP_3189_elements(258)); -- 
    cr_5339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(258), ack => RPIPE_input_done_pipe_2274_inst_req_1); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/RPIPE_input_done_pipe_2274_update_completed_
      -- 
    ca_5340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2274_inst_ack_1, ack => convolution3D_CP_3189_elements(259)); -- 
    -- CP-element group 260:  join  transition  place  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	257 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (7) 
      -- CP-element group 260: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275__exit__
      -- CP-element group 260: 	 branch_block_stmt_1049/assign_stmt_2279__entry__
      -- CP-element group 260: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_1049/assign_stmt_2279/$entry
      -- CP-element group 260: 	 branch_block_stmt_1049/assign_stmt_2272_to_assign_stmt_2275/$exit
      -- 
    rr_5351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(260), ack => RPIPE_input_done_pipe_2278_inst_req_0); -- 
    convolution3D_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(257) & convolution3D_CP_3189_elements(259);
      gj_convolution3D_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Sample/ra
      -- CP-element group 261: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_update_start_
      -- CP-element group 261: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_sample_completed_
      -- 
    ra_5352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2278_inst_ack_0, ack => convolution3D_CP_3189_elements(261)); -- 
    cr_5356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(261), ack => RPIPE_input_done_pipe_2278_inst_req_1); -- 
    -- CP-element group 262:  fork  transition  place  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	273 
    -- CP-element group 262: 	269 
    -- CP-element group 262: 	270 
    -- CP-element group 262: 	266 
    -- CP-element group 262: 	267 
    -- CP-element group 262: 	268 
    -- CP-element group 262: 	263 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (31) 
      -- CP-element group 262: 	 branch_block_stmt_1049/assign_stmt_2279__exit__
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327__entry__
      -- CP-element group 262: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_Update/ca
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Sample/crr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/assign_stmt_2279/RPIPE_input_done_pipe_2278_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/assign_stmt_2279/$exit
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Update/ccr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Update/ccr
      -- CP-element group 262: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Update/$entry
      -- 
    ca_5357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2278_inst_ack_1, ack => convolution3D_CP_3189_elements(262)); -- 
    crr_5368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => call_stmt_2282_call_req_0); -- 
    cr_5415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => type_cast_2299_inst_req_1); -- 
    rr_5410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => type_cast_2299_inst_req_0); -- 
    cr_5401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => type_cast_2295_inst_req_1); -- 
    rr_5396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => type_cast_2295_inst_req_0); -- 
    cr_5387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => type_cast_2286_inst_req_1); -- 
    ccr_5429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => call_stmt_2327_call_req_1); -- 
    ccr_5373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(262), ack => call_stmt_2282_call_req_1); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Sample/cra
      -- 
    cra_5369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2282_call_ack_0, ack => convolution3D_CP_3189_elements(263)); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Sample/rr
      -- CP-element group 264: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Update/cca
      -- CP-element group 264: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2282_Update/$exit
      -- 
    cca_5374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2282_call_ack_1, ack => convolution3D_CP_3189_elements(264)); -- 
    rr_5382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(264), ack => type_cast_2286_inst_req_0); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Sample/ra
      -- CP-element group 265: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_sample_completed_
      -- 
    ra_5383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2286_inst_ack_0, ack => convolution3D_CP_3189_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	262 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	274 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Update/ca
      -- CP-element group 266: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2286_update_completed_
      -- 
    ca_5388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2286_inst_ack_1, ack => convolution3D_CP_3189_elements(266)); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	262 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Sample/ra
      -- CP-element group 267: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_sample_completed_
      -- 
    ra_5397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_0, ack => convolution3D_CP_3189_elements(267)); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	262 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	271 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2295_update_completed_
      -- 
    ca_5402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_1, ack => convolution3D_CP_3189_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	262 
    -- CP-element group 269: successors 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Sample/ra
      -- CP-element group 269: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_sample_completed_
      -- 
    ra_5411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2299_inst_ack_0, ack => convolution3D_CP_3189_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	262 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Update/ca
      -- CP-element group 270: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/type_cast_2299_update_completed_
      -- 
    ca_5416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2299_inst_ack_1, ack => convolution3D_CP_3189_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: 	268 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Sample/crr
      -- 
    crr_5424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(271), ack => call_stmt_2327_call_req_0); -- 
    convolution3D_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(270) & convolution3D_CP_3189_elements(268);
      gj_convolution3D_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Sample/cra
      -- 
    cra_5425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2327_call_ack_0, ack => convolution3D_CP_3189_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	262 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Update/cca
      -- CP-element group 273: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/call_stmt_2327_Update/$exit
      -- 
    cca_5430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2327_call_ack_1, ack => convolution3D_CP_3189_elements(273)); -- 
    -- CP-element group 274:  join  fork  transition  place  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: 	266 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274: 	276 
    -- CP-element group 274: 	289 
    -- CP-element group 274: 	290 
    -- CP-element group 274: 	285 
    -- CP-element group 274: 	286 
    -- CP-element group 274: 	287 
    -- CP-element group 274: 	288 
    -- CP-element group 274: 	277 
    -- CP-element group 274: 	278 
    -- CP-element group 274: 	279 
    -- CP-element group 274: 	280 
    -- CP-element group 274: 	281 
    -- CP-element group 274: 	282 
    -- CP-element group 274: 	283 
    -- CP-element group 274: 	284 
    -- CP-element group 274:  members (52) 
      -- CP-element group 274: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327__exit__
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426__entry__
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/call_stmt_2282_to_call_stmt_2327/$exit
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Sample/rr
      -- 
    cr_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2371_inst_req_1); -- 
    cr_5474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2351_inst_req_1); -- 
    rr_5455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2341_inst_req_0); -- 
    rr_5539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2401_inst_req_0); -- 
    cr_5446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2331_inst_req_1); -- 
    cr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2391_inst_req_1); -- 
    rr_5497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2371_inst_req_0); -- 
    cr_5544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2401_inst_req_1); -- 
    rr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2391_inst_req_0); -- 
    rr_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2331_inst_req_0); -- 
    rr_5469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2351_inst_req_0); -- 
    cr_5516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2381_inst_req_1); -- 
    cr_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2361_inst_req_1); -- 
    cr_5460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2341_inst_req_1); -- 
    rr_5511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2381_inst_req_0); -- 
    rr_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(274), ack => type_cast_2361_inst_req_0); -- 
    convolution3D_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(273) & convolution3D_CP_3189_elements(266);
      gj_convolution3D_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Sample/ra
      -- CP-element group 275: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_sample_completed_
      -- 
    ra_5442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_0, ack => convolution3D_CP_3189_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	311 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Update/ca
      -- CP-element group 276: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2331_update_completed_
      -- 
    ca_5447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_1, ack => convolution3D_CP_3189_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	274 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Sample/ra
      -- 
    ra_5456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_0, ack => convolution3D_CP_3189_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	274 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	308 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Update/ca
      -- CP-element group 278: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2341_Update/$exit
      -- 
    ca_5461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_1, ack => convolution3D_CP_3189_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	274 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_sample_completed_
      -- 
    ra_5470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_0, ack => convolution3D_CP_3189_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	274 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	305 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_Update/ca
      -- CP-element group 280: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2351_update_completed_
      -- 
    ca_5475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_1, ack => convolution3D_CP_3189_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	274 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Sample/$exit
      -- 
    ra_5484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2361_inst_ack_0, ack => convolution3D_CP_3189_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	274 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	302 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2361_Update/$exit
      -- 
    ca_5489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2361_inst_ack_1, ack => convolution3D_CP_3189_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	274 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Sample/ra
      -- CP-element group 283: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_sample_completed_
      -- 
    ra_5498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_0, ack => convolution3D_CP_3189_elements(283)); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	274 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	299 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Update/ca
      -- CP-element group 284: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2371_update_completed_
      -- 
    ca_5503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_1, ack => convolution3D_CP_3189_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	274 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Sample/ra
      -- CP-element group 285: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Sample/$exit
      -- 
    ra_5512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2381_inst_ack_0, ack => convolution3D_CP_3189_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	274 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	296 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Update/ca
      -- CP-element group 286: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2381_Update/$exit
      -- 
    ca_5517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2381_inst_ack_1, ack => convolution3D_CP_3189_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	274 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Sample/ra
      -- CP-element group 287: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_sample_completed_
      -- 
    ra_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2391_inst_ack_0, ack => convolution3D_CP_3189_elements(287)); -- 
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	274 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	293 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Update/ca
      -- CP-element group 288: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2391_update_completed_
      -- 
    ca_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2391_inst_ack_1, ack => convolution3D_CP_3189_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	274 
    -- CP-element group 289: successors 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Sample/ra
      -- CP-element group 289: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_sample_completed_
      -- 
    ra_5540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_0, ack => convolution3D_CP_3189_elements(289)); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	274 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/type_cast_2401_Update/ca
      -- CP-element group 290: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Sample/req
      -- 
    ca_5545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_1, ack => convolution3D_CP_3189_elements(290)); -- 
    req_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(290), ack => WPIPE_maxpool_output_pipe_2403_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_update_start_
      -- CP-element group 291: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Update/req
      -- 
    ack_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2403_inst_ack_0, ack => convolution3D_CP_3189_elements(291)); -- 
    req_5558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(291), ack => WPIPE_maxpool_output_pipe_2403_inst_req_1); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2403_Update/ack
      -- 
    ack_5559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2403_inst_ack_1, ack => convolution3D_CP_3189_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: 	288 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Sample/req
      -- 
    req_5567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(293), ack => WPIPE_maxpool_output_pipe_2406_inst_req_0); -- 
    convolution3D_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(292) & convolution3D_CP_3189_elements(288);
      gj_convolution3D_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_sample_completed_
      -- CP-element group 294: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_update_start_
      -- CP-element group 294: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Sample/ack
      -- CP-element group 294: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Update/req
      -- 
    ack_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2406_inst_ack_0, ack => convolution3D_CP_3189_elements(294)); -- 
    req_5572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(294), ack => WPIPE_maxpool_output_pipe_2406_inst_req_1); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_update_completed_
      -- CP-element group 295: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2406_Update/ack
      -- 
    ack_5573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2406_inst_ack_1, ack => convolution3D_CP_3189_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: 	286 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Sample/req
      -- 
    req_5581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(296), ack => WPIPE_maxpool_output_pipe_2409_inst_req_0); -- 
    convolution3D_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(295) & convolution3D_CP_3189_elements(286);
      gj_convolution3D_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_update_start_
      -- CP-element group 297: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Update/req
      -- 
    ack_5582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2409_inst_ack_0, ack => convolution3D_CP_3189_elements(297)); -- 
    req_5586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(297), ack => WPIPE_maxpool_output_pipe_2409_inst_req_1); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2409_Update/ack
      -- 
    ack_5587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2409_inst_ack_1, ack => convolution3D_CP_3189_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	284 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_sample_start_
      -- CP-element group 299: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Sample/req
      -- 
    req_5595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(299), ack => WPIPE_maxpool_output_pipe_2412_inst_req_0); -- 
    convolution3D_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(284) & convolution3D_CP_3189_elements(298);
      gj_convolution3D_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_update_start_
      -- CP-element group 300: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Sample/ack
      -- CP-element group 300: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Update/req
      -- 
    ack_5596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2412_inst_ack_0, ack => convolution3D_CP_3189_elements(300)); -- 
    req_5600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(300), ack => WPIPE_maxpool_output_pipe_2412_inst_req_1); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2412_Update/ack
      -- 
    ack_5601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2412_inst_ack_1, ack => convolution3D_CP_3189_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	282 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Sample/req
      -- 
    req_5609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(302), ack => WPIPE_maxpool_output_pipe_2415_inst_req_0); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(282) & convolution3D_CP_3189_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_update_start_
      -- CP-element group 303: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Update/req
      -- 
    ack_5610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2415_inst_ack_0, ack => convolution3D_CP_3189_elements(303)); -- 
    req_5614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(303), ack => WPIPE_maxpool_output_pipe_2415_inst_req_1); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2415_Update/ack
      -- 
    ack_5615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2415_inst_ack_1, ack => convolution3D_CP_3189_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	280 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Sample/req
      -- 
    req_5623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(305), ack => WPIPE_maxpool_output_pipe_2418_inst_req_0); -- 
    convolution3D_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(280) & convolution3D_CP_3189_elements(304);
      gj_convolution3D_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_update_start_
      -- CP-element group 306: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Sample/ack
      -- CP-element group 306: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Update/req
      -- 
    ack_5624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2418_inst_ack_0, ack => convolution3D_CP_3189_elements(306)); -- 
    req_5628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(306), ack => WPIPE_maxpool_output_pipe_2418_inst_req_1); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2418_Update/ack
      -- 
    ack_5629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2418_inst_ack_1, ack => convolution3D_CP_3189_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	278 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Sample/req
      -- 
    req_5637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(308), ack => WPIPE_maxpool_output_pipe_2421_inst_req_0); -- 
    convolution3D_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(278) & convolution3D_CP_3189_elements(307);
      gj_convolution3D_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_update_start_
      -- CP-element group 309: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Update/req
      -- 
    ack_5638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2421_inst_ack_0, ack => convolution3D_CP_3189_elements(309)); -- 
    req_5642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(309), ack => WPIPE_maxpool_output_pipe_2421_inst_req_1); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2421_Update/ack
      -- 
    ack_5643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2421_inst_ack_1, ack => convolution3D_CP_3189_elements(310)); -- 
    -- CP-element group 311:  join  transition  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	276 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_sample_start_
      -- CP-element group 311: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Sample/req
      -- 
    req_5651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(311), ack => WPIPE_maxpool_output_pipe_2424_inst_req_0); -- 
    convolution3D_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(276) & convolution3D_CP_3189_elements(310);
      gj_convolution3D_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_update_start_
      -- CP-element group 312: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Sample/ack
      -- CP-element group 312: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Update/req
      -- 
    ack_5652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2424_inst_ack_0, ack => convolution3D_CP_3189_elements(312)); -- 
    req_5656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(312), ack => WPIPE_maxpool_output_pipe_2424_inst_req_1); -- 
    -- CP-element group 313:  transition  place  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (16) 
      -- CP-element group 313: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426__exit__
      -- CP-element group 313: 	 branch_block_stmt_1049/return__
      -- CP-element group 313: 	 branch_block_stmt_1049/merge_stmt_2428__exit__
      -- CP-element group 313: 	 $exit
      -- CP-element group 313: 	 branch_block_stmt_1049/$exit
      -- CP-element group 313: 	 branch_block_stmt_1049/branch_block_stmt_1049__exit__
      -- CP-element group 313: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/$exit
      -- CP-element group 313: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_1049/assign_stmt_2332_to_assign_stmt_2426/WPIPE_maxpool_output_pipe_2424_Update/ack
      -- CP-element group 313: 	 branch_block_stmt_1049/return___PhiReq/$entry
      -- CP-element group 313: 	 branch_block_stmt_1049/return___PhiReq/$exit
      -- CP-element group 313: 	 branch_block_stmt_1049/merge_stmt_2428_PhiReqMerge
      -- CP-element group 313: 	 branch_block_stmt_1049/merge_stmt_2428_PhiAck/$entry
      -- CP-element group 313: 	 branch_block_stmt_1049/merge_stmt_2428_PhiAck/$exit
      -- CP-element group 313: 	 branch_block_stmt_1049/merge_stmt_2428_PhiAck/dummy
      -- 
    ack_5657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2424_inst_ack_1, ack => convolution3D_CP_3189_elements(313)); -- 
    -- CP-element group 314:  transition  output  delay-element  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	86 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	318 
    -- CP-element group 314:  members (5) 
      -- CP-element group 314: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/$exit
      -- CP-element group 314: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1358/$exit
      -- CP-element group 314: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/$exit
      -- CP-element group 314: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1362_konst_delay_trans
      -- CP-element group 314: 	 branch_block_stmt_1049/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_req
      -- 
    phi_stmt_1358_req_5680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1358_req_5680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(314), ack => phi_stmt_1358_req_0); -- 
    -- Element group convolution3D_CP_3189_elements(314) is a control-delay.
    cp_element_314_delay: control_delay_element  generic map(name => " 314_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(86), ack => convolution3D_CP_3189_elements(314), clk => clk, reset =>reset);
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	128 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Sample/ra
      -- 
    ra_5700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1364_inst_ack_0, ack => convolution3D_CP_3189_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	128 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/Update/ca
      -- 
    ca_5705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1364_inst_ack_1, ack => convolution3D_CP_3189_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 317: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/$exit
      -- CP-element group 317: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/$exit
      -- CP-element group 317: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/$exit
      -- CP-element group 317: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_sources/type_cast_1364/SplitProtocol/$exit
      -- CP-element group 317: 	 branch_block_stmt_1049/forx_xbody_forx_xbody_PhiReq/phi_stmt_1358/phi_stmt_1358_req
      -- 
    phi_stmt_1358_req_5706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1358_req_5706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(317), ack => phi_stmt_1358_req_1); -- 
    convolution3D_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(315) & convolution3D_CP_3189_elements(316);
      gj_convolution3D_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  merge  transition  place  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	314 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_1049/merge_stmt_1357_PhiReqMerge
      -- CP-element group 318: 	 branch_block_stmt_1049/merge_stmt_1357_PhiAck/$entry
      -- 
    convolution3D_CP_3189_elements(318) <= OrReduce(convolution3D_CP_3189_elements(314) & convolution3D_CP_3189_elements(317));
    -- CP-element group 319:  fork  transition  place  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	110 
    -- CP-element group 319: 	122 
    -- CP-element group 319: 	114 
    -- CP-element group 319: 	125 
    -- CP-element group 319: 	118 
    -- CP-element group 319: 	87 
    -- CP-element group 319: 	88 
    -- CP-element group 319: 	90 
    -- CP-element group 319: 	91 
    -- CP-element group 319: 	94 
    -- CP-element group 319: 	98 
    -- CP-element group 319: 	102 
    -- CP-element group 319: 	106 
    -- CP-element group 319:  members (56) 
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1481_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/merge_stmt_1357__exit__
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520__entry__
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_resized_1
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_scaled_1
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_computed_1
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1463_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_resize_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_resize_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_resize_1/index_resize_req
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_resize_1/index_resize_ack
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_scale_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_scale_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_scale_1/scale_rename_req
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_index_scale_1/scale_rename_ack
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_update_start
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Sample/req
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/array_obj_ref_1370_final_index_sum_regn_Update/req
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/word_access_complete/word_0/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_complete/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/addr_of_1371_complete/req
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/word_access_complete/word_0/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_sample_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/RPIPE_maxpool_input_pipe_1374_Sample/rr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/word_access_complete/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1378_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/ptr_deref_1507_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1499_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1391_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1409_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1427_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1049/assign_stmt_1372_to_assign_stmt_1520/type_cast_1445_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1049/merge_stmt_1357_PhiAck/$exit
      -- CP-element group 319: 	 branch_block_stmt_1049/merge_stmt_1357_PhiAck/phi_stmt_1358_ack
      -- 
    phi_stmt_1358_ack_5711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1358_ack_0, ack => convolution3D_CP_3189_elements(319)); -- 
    cr_4087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1463_inst_req_1); -- 
    cr_4115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1481_inst_req_1); -- 
    cr_4143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1499_inst_req_1); -- 
    req_3899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => array_obj_ref_1370_index_offset_req_0); -- 
    req_3904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => array_obj_ref_1370_index_offset_req_1); -- 
    cr_4193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => ptr_deref_1507_store_0_req_1); -- 
    req_3919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => addr_of_1371_final_reg_req_1); -- 
    rr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => RPIPE_maxpool_input_pipe_1374_inst_req_0); -- 
    cr_3947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1378_inst_req_1); -- 
    cr_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1391_inst_req_1); -- 
    cr_4003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1409_inst_req_1); -- 
    cr_4031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1427_inst_req_1); -- 
    cr_4059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(319), ack => type_cast_1445_inst_req_1); -- 
    -- CP-element group 320:  transition  output  delay-element  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	76 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	324 
    -- CP-element group 320:  members (5) 
      -- CP-element group 320: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/$exit
      -- CP-element group 320: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/phi_stmt_1552/$exit
      -- CP-element group 320: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$exit
      -- CP-element group 320: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558_konst_delay_trans
      -- CP-element group 320: 	 branch_block_stmt_1049/entry_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_req
      -- 
    phi_stmt_1552_req_5734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1552_req_5734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(320), ack => phi_stmt_1552_req_1); -- 
    -- Element group convolution3D_CP_3189_elements(320) is a control-delay.
    cp_element_320_delay: control_delay_element  generic map(name => " 320_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(76), ack => convolution3D_CP_3189_elements(320), clk => clk, reset =>reset);
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	127 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Sample/ra
      -- 
    ra_5754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1555_inst_ack_0, ack => convolution3D_CP_3189_elements(321)); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	127 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/Update/ca
      -- 
    ca_5759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1555_inst_ack_1, ack => convolution3D_CP_3189_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 323: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/$exit
      -- CP-element group 323: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$exit
      -- CP-element group 323: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/$exit
      -- CP-element group 323: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1555/SplitProtocol/$exit
      -- CP-element group 323: 	 branch_block_stmt_1049/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1552/phi_stmt_1552_req
      -- 
    phi_stmt_1552_req_5760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1552_req_5760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(323), ack => phi_stmt_1552_req_0); -- 
    convolution3D_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(321) & convolution3D_CP_3189_elements(322);
      gj_convolution3D_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  merge  transition  place  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	320 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (2) 
      -- CP-element group 324: 	 branch_block_stmt_1049/merge_stmt_1551_PhiReqMerge
      -- CP-element group 324: 	 branch_block_stmt_1049/merge_stmt_1551_PhiAck/$entry
      -- 
    convolution3D_CP_3189_elements(324) <= OrReduce(convolution3D_CP_3189_elements(320) & convolution3D_CP_3189_elements(323));
    -- CP-element group 325:  branch  transition  place  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	129 
    -- CP-element group 325: 	130 
    -- CP-element group 325:  members (15) 
      -- CP-element group 325: 	 branch_block_stmt_1049/merge_stmt_1551__exit__
      -- CP-element group 325: 	 branch_block_stmt_1049/assign_stmt_1565_to_assign_stmt_1571__entry__
      -- CP-element group 325: 	 branch_block_stmt_1049/assign_stmt_1565_to_assign_stmt_1571__exit__
      -- CP-element group 325: 	 branch_block_stmt_1049/if_stmt_1572__entry__
      -- CP-element group 325: 	 branch_block_stmt_1049/if_stmt_1572_else_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_1049/if_stmt_1572_if_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_1049/if_stmt_1572_eval_test/branch_req
      -- CP-element group 325: 	 branch_block_stmt_1049/if_stmt_1572_eval_test/$exit
      -- CP-element group 325: 	 branch_block_stmt_1049/if_stmt_1572_eval_test/$entry
      -- CP-element group 325: 	 branch_block_stmt_1049/if_stmt_1572_dead_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_1049/assign_stmt_1565_to_assign_stmt_1571/$exit
      -- CP-element group 325: 	 branch_block_stmt_1049/assign_stmt_1565_to_assign_stmt_1571/$entry
      -- CP-element group 325: 	 branch_block_stmt_1049/R_tobool_1573_place
      -- CP-element group 325: 	 branch_block_stmt_1049/merge_stmt_1551_PhiAck/$exit
      -- CP-element group 325: 	 branch_block_stmt_1049/merge_stmt_1551_PhiAck/phi_stmt_1552_ack
      -- 
    phi_stmt_1552_ack_5765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1552_ack_0, ack => convolution3D_CP_3189_elements(325)); -- 
    branch_req_4227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(325), ack => if_stmt_1572_branch_req_0); -- 
    -- CP-element group 326:  transition  output  delay-element  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	130 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (4) 
      -- CP-element group 326: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/$exit
      -- CP-element group 326: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/$exit
      -- CP-element group 326: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1597_konst_delay_trans
      -- CP-element group 326: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_req
      -- 
    phi_stmt_1593_req_5788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1593_req_5788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(326), ack => phi_stmt_1593_req_0); -- 
    -- Element group convolution3D_CP_3189_elements(326) is a control-delay.
    cp_element_326_delay: control_delay_element  generic map(name => " 326_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(130), ack => convolution3D_CP_3189_elements(326), clk => clk, reset =>reset);
    -- CP-element group 327:  transition  output  delay-element  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	130 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (4) 
      -- CP-element group 327: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/$exit
      -- CP-element group 327: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$exit
      -- CP-element group 327: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1604_konst_delay_trans
      -- CP-element group 327: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_req
      -- 
    phi_stmt_1600_req_5796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1600_req_5796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(327), ack => phi_stmt_1600_req_0); -- 
    -- Element group convolution3D_CP_3189_elements(327) is a control-delay.
    cp_element_327_delay: control_delay_element  generic map(name => " 327_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(130), ack => convolution3D_CP_3189_elements(327), clk => clk, reset =>reset);
    -- CP-element group 328:  join  transition  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	336 
    -- CP-element group 328:  members (1) 
      -- CP-element group 328: 	 branch_block_stmt_1049/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(326) & convolution3D_CP_3189_elements(327);
      gj_convolution3D_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	138 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (2) 
      -- CP-element group 329: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Sample/ra
      -- 
    ra_5816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1599_inst_ack_0, ack => convolution3D_CP_3189_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	138 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (2) 
      -- CP-element group 330: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/Update/ca
      -- 
    ca_5821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1599_inst_ack_1, ack => convolution3D_CP_3189_elements(330)); -- 
    -- CP-element group 331:  join  transition  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	335 
    -- CP-element group 331:  members (5) 
      -- CP-element group 331: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/$exit
      -- CP-element group 331: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/$exit
      -- CP-element group 331: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/$exit
      -- CP-element group 331: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_sources/type_cast_1599/SplitProtocol/$exit
      -- CP-element group 331: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1593/phi_stmt_1593_req
      -- 
    phi_stmt_1593_req_5822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1593_req_5822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(331), ack => phi_stmt_1593_req_1); -- 
    convolution3D_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(329) & convolution3D_CP_3189_elements(330);
      gj_convolution3D_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	138 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	334 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/ra
      -- 
    ra_5839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_0, ack => convolution3D_CP_3189_elements(332)); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	138 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (2) 
      -- CP-element group 333: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/ca
      -- 
    ca_5844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_1, ack => convolution3D_CP_3189_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	332 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (5) 
      -- CP-element group 334: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/$exit
      -- CP-element group 334: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$exit
      -- CP-element group 334: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/$exit
      -- CP-element group 334: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/$exit
      -- CP-element group 334: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1600/phi_stmt_1600_req
      -- 
    phi_stmt_1600_req_5845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1600_req_5845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(334), ack => phi_stmt_1600_req_1); -- 
    convolution3D_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(332) & convolution3D_CP_3189_elements(333);
      gj_convolution3D_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	331 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (1) 
      -- CP-element group 335: 	 branch_block_stmt_1049/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(331) & convolution3D_CP_3189_elements(334);
      gj_convolution3D_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  merge  fork  transition  place  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	328 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336: 	338 
    -- CP-element group 336:  members (2) 
      -- CP-element group 336: 	 branch_block_stmt_1049/merge_stmt_1592_PhiReqMerge
      -- CP-element group 336: 	 branch_block_stmt_1049/merge_stmt_1592_PhiAck/$entry
      -- 
    convolution3D_CP_3189_elements(336) <= OrReduce(convolution3D_CP_3189_elements(328) & convolution3D_CP_3189_elements(335));
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337:  members (1) 
      -- CP-element group 337: 	 branch_block_stmt_1049/merge_stmt_1592_PhiAck/phi_stmt_1593_ack
      -- 
    phi_stmt_1593_ack_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1593_ack_0, ack => convolution3D_CP_3189_elements(337)); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (1) 
      -- CP-element group 338: 	 branch_block_stmt_1049/merge_stmt_1592_PhiAck/phi_stmt_1600_ack
      -- 
    phi_stmt_1600_ack_5851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1600_ack_0, ack => convolution3D_CP_3189_elements(338)); -- 
    -- CP-element group 339:  join  fork  transition  place  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	131 
    -- CP-element group 339: 	134 
    -- CP-element group 339: 	135 
    -- CP-element group 339: 	136 
    -- CP-element group 339:  members (16) 
      -- CP-element group 339: 	 branch_block_stmt_1049/merge_stmt_1592__exit__
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646__entry__
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/$entry
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Update/cr
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Sample/rr
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_update_start_
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1640_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Update/cr
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/type_cast_1625_update_start_
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Sample/rr
      -- CP-element group 339: 	 branch_block_stmt_1049/assign_stmt_1613_to_assign_stmt_1646/RPIPE_maxpool_input_pipe_1621_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_1049/merge_stmt_1592_PhiAck/$exit
      -- 
    cr_4285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(339), ack => type_cast_1640_inst_req_1); -- 
    rr_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(339), ack => type_cast_1640_inst_req_0); -- 
    cr_4271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(339), ack => type_cast_1625_inst_req_1); -- 
    rr_4252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(339), ack => RPIPE_maxpool_input_pipe_1621_inst_req_0); -- 
    convolution3D_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(337) & convolution3D_CP_3189_elements(338);
      gj_convolution3D_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	139 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (2) 
      -- CP-element group 340: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Sample/ra
      -- 
    ra_5875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1657_inst_ack_0, ack => convolution3D_CP_3189_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	139 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (2) 
      -- CP-element group 341: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/Update/ca
      -- 
    ca_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1657_inst_ack_1, ack => convolution3D_CP_3189_elements(341)); -- 
    -- CP-element group 342:  join  transition  place  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (8) 
      -- CP-element group 342: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 342: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/$exit
      -- CP-element group 342: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/$exit
      -- CP-element group 342: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/$exit
      -- CP-element group 342: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_sources/type_cast_1657/SplitProtocol/$exit
      -- CP-element group 342: 	 branch_block_stmt_1049/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1654/phi_stmt_1654_req
      -- CP-element group 342: 	 branch_block_stmt_1049/merge_stmt_1653_PhiReqMerge
      -- CP-element group 342: 	 branch_block_stmt_1049/merge_stmt_1653_PhiAck/$entry
      -- 
    phi_stmt_1654_req_5881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1654_req_5881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(342), ack => phi_stmt_1654_req_0); -- 
    convolution3D_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(340) & convolution3D_CP_3189_elements(341);
      gj_convolution3D_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	140 
    -- CP-element group 343: 	141 
    -- CP-element group 343: 	143 
    -- CP-element group 343: 	145 
    -- CP-element group 343:  members (29) 
      -- CP-element group 343: 	 branch_block_stmt_1049/merge_stmt_1653__exit__
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_resize_1/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692__entry__
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_computed_1
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_scale_1/scale_rename_ack
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/word_access_complete/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_resized_1
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_scaled_1
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_update_start_
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_update_start_
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_scale_1/scale_rename_req
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_complete/req
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_scale_1/$exit
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/addr_of_1687_complete/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/word_access_complete/word_0/cr
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_scale_1/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_resize_1/index_resize_ack
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_resize_1/index_resize_req
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Update/req
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/ptr_deref_1690_Update/word_access_complete/word_0/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Sample/req
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_index_resize_1/$exit
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_1049/assign_stmt_1664_to_assign_stmt_1692/array_obj_ref_1686_final_index_sum_regn_update_start
      -- CP-element group 343: 	 branch_block_stmt_1049/merge_stmt_1653_PhiAck/$exit
      -- CP-element group 343: 	 branch_block_stmt_1049/merge_stmt_1653_PhiAck/phi_stmt_1654_ack
      -- 
    phi_stmt_1654_ack_5886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1654_ack_0, ack => convolution3D_CP_3189_elements(343)); -- 
    req_4353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(343), ack => addr_of_1687_final_reg_req_1); -- 
    cr_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(343), ack => ptr_deref_1690_store_0_req_1); -- 
    req_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(343), ack => array_obj_ref_1686_index_offset_req_1); -- 
    req_4333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(343), ack => array_obj_ref_1686_index_offset_req_0); -- 
    -- CP-element group 344:  merge  fork  transition  place  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	129 
    -- CP-element group 344: 	146 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	150 
    -- CP-element group 344: 	151 
    -- CP-element group 344: 	152 
    -- CP-element group 344: 	147 
    -- CP-element group 344: 	148 
    -- CP-element group 344: 	149 
    -- CP-element group 344:  members (25) 
      -- CP-element group 344: 	 branch_block_stmt_1049/merge_stmt_1694__exit__
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742__entry__
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Update/cr
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_update_start_
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Update/cr
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Sample/rr
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Update/cr
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_update_start_
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1697_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Sample/rr
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1705_Sample/rr
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_update_start_
      -- CP-element group 344: 	 branch_block_stmt_1049/assign_stmt_1698_to_assign_stmt_1742/type_cast_1701_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/merge_stmt_1694_PhiReqMerge
      -- CP-element group 344: 	 branch_block_stmt_1049/merge_stmt_1694_PhiAck/$entry
      -- CP-element group 344: 	 branch_block_stmt_1049/merge_stmt_1694_PhiAck/$exit
      -- CP-element group 344: 	 branch_block_stmt_1049/merge_stmt_1694_PhiAck/dummy
      -- 
    cr_4448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(344), ack => type_cast_1705_inst_req_1); -- 
    cr_4420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(344), ack => type_cast_1697_inst_req_1); -- 
    rr_4415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(344), ack => type_cast_1697_inst_req_0); -- 
    cr_4434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(344), ack => type_cast_1701_inst_req_1); -- 
    rr_4429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(344), ack => type_cast_1701_inst_req_0); -- 
    rr_4443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(344), ack => type_cast_1705_inst_req_0); -- 
    convolution3D_CP_3189_elements(344) <= OrReduce(convolution3D_CP_3189_elements(129) & convolution3D_CP_3189_elements(146));
    -- CP-element group 345:  transition  output  delay-element  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	166 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	349 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- CP-element group 345: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1819/$exit
      -- CP-element group 345: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$exit
      -- CP-element group 345: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825_konst_delay_trans
      -- CP-element group 345: 	 branch_block_stmt_1049/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_req
      -- 
    phi_stmt_1819_req_5920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1819_req_5920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(345), ack => phi_stmt_1819_req_1); -- 
    -- Element group convolution3D_CP_3189_elements(345) is a control-delay.
    cp_element_345_delay: control_delay_element  generic map(name => " 345_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(166), ack => convolution3D_CP_3189_elements(345), clk => clk, reset =>reset);
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	208 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Sample/ra
      -- 
    ra_5940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_0, ack => convolution3D_CP_3189_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	208 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (2) 
      -- CP-element group 347: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/Update/ca
      -- 
    ca_5945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_1, ack => convolution3D_CP_3189_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (6) 
      -- CP-element group 348: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 348: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/$exit
      -- CP-element group 348: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$exit
      -- CP-element group 348: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/$exit
      -- CP-element group 348: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1822/SplitProtocol/$exit
      -- CP-element group 348: 	 branch_block_stmt_1049/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1819/phi_stmt_1819_req
      -- 
    phi_stmt_1819_req_5946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1819_req_5946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(348), ack => phi_stmt_1819_req_0); -- 
    convolution3D_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(346) & convolution3D_CP_3189_elements(347);
      gj_convolution3D_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  merge  transition  place  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	345 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (2) 
      -- CP-element group 349: 	 branch_block_stmt_1049/merge_stmt_1818_PhiReqMerge
      -- CP-element group 349: 	 branch_block_stmt_1049/merge_stmt_1818_PhiAck/$entry
      -- 
    convolution3D_CP_3189_elements(349) <= OrReduce(convolution3D_CP_3189_elements(345) & convolution3D_CP_3189_elements(348));
    -- CP-element group 350:  fork  transition  place  input  output  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	174 
    -- CP-element group 350: 	178 
    -- CP-element group 350: 	167 
    -- CP-element group 350: 	168 
    -- CP-element group 350: 	186 
    -- CP-element group 350: 	170 
    -- CP-element group 350: 	171 
    -- CP-element group 350: 	190 
    -- CP-element group 350: 	198 
    -- CP-element group 350: 	182 
    -- CP-element group 350: 	205 
    -- CP-element group 350: 	194 
    -- CP-element group 350: 	202 
    -- CP-element group 350:  members (56) 
      -- CP-element group 350: 	 branch_block_stmt_1049/merge_stmt_1818__exit__
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981__entry__
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_resized_1
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_scaled_1
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_computed_1
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_resize_1/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_resize_1/$exit
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_resize_1/index_resize_req
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_resize_1/index_resize_ack
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_scale_1/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_scale_1/$exit
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_scale_1/scale_rename_req
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_index_scale_1/scale_rename_ack
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_update_start
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Sample/req
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/array_obj_ref_1831_final_index_sum_regn_Update/req
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/addr_of_1832_complete/req
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_sample_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/RPIPE_maxpool_input_pipe_1835_Sample/rr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1839_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1852_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1870_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1888_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1906_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1924_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1942_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/type_cast_1960_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/word_access_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/word_access_complete/word_0/$entry
      -- CP-element group 350: 	 branch_block_stmt_1049/assign_stmt_1833_to_assign_stmt_1981/ptr_deref_1968_Update/word_access_complete/word_0/cr
      -- CP-element group 350: 	 branch_block_stmt_1049/merge_stmt_1818_PhiAck/$exit
      -- CP-element group 350: 	 branch_block_stmt_1049/merge_stmt_1818_PhiAck/phi_stmt_1819_ack
      -- 
    phi_stmt_1819_ack_5951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1819_ack_0, ack => convolution3D_CP_3189_elements(350)); -- 
    req_4569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => array_obj_ref_1831_index_offset_req_0); -- 
    req_4574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => array_obj_ref_1831_index_offset_req_1); -- 
    req_4589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => addr_of_1832_final_reg_req_1); -- 
    rr_4598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => RPIPE_maxpool_input_pipe_1835_inst_req_0); -- 
    cr_4617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1839_inst_req_1); -- 
    cr_4645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1852_inst_req_1); -- 
    cr_4673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1870_inst_req_1); -- 
    cr_4701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1888_inst_req_1); -- 
    cr_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1906_inst_req_1); -- 
    cr_4757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1924_inst_req_1); -- 
    cr_4785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1942_inst_req_1); -- 
    cr_4813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => type_cast_1960_inst_req_1); -- 
    cr_4863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(350), ack => ptr_deref_1968_store_0_req_1); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	207 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (2) 
      -- CP-element group 351: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Sample/ra
      -- 
    ra_5983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2016_inst_ack_0, ack => convolution3D_CP_3189_elements(351)); -- 
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	207 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (2) 
      -- CP-element group 352: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/Update/ca
      -- 
    ca_5988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2016_inst_ack_1, ack => convolution3D_CP_3189_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (6) 
      -- CP-element group 353: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- CP-element group 353: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/$exit
      -- CP-element group 353: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/$exit
      -- CP-element group 353: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/$exit
      -- CP-element group 353: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2016/SplitProtocol/$exit
      -- CP-element group 353: 	 branch_block_stmt_1049/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_req
      -- 
    phi_stmt_2013_req_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2013_req_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(353), ack => phi_stmt_2013_req_0); -- 
    convolution3D_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(351) & convolution3D_CP_3189_elements(352);
      gj_convolution3D_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  transition  output  delay-element  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	155 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (5) 
      -- CP-element group 354: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/$exit
      -- CP-element group 354: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/phi_stmt_2013/$exit
      -- CP-element group 354: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/$exit
      -- CP-element group 354: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_sources/type_cast_2019_konst_delay_trans
      -- CP-element group 354: 	 branch_block_stmt_1049/ifx_xend_forx_xend215_PhiReq/phi_stmt_2013/phi_stmt_2013_req
      -- 
    phi_stmt_2013_req_6000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2013_req_6000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(354), ack => phi_stmt_2013_req_1); -- 
    -- Element group convolution3D_CP_3189_elements(354) is a control-delay.
    cp_element_354_delay: control_delay_element  generic map(name => " 354_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(155), ack => convolution3D_CP_3189_elements(354), clk => clk, reset =>reset);
    -- CP-element group 355:  merge  transition  place  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (2) 
      -- CP-element group 355: 	 branch_block_stmt_1049/merge_stmt_2012_PhiReqMerge
      -- CP-element group 355: 	 branch_block_stmt_1049/merge_stmt_2012_PhiAck/$entry
      -- 
    convolution3D_CP_3189_elements(355) <= OrReduce(convolution3D_CP_3189_elements(353) & convolution3D_CP_3189_elements(354));
    -- CP-element group 356:  branch  transition  place  input  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	209 
    -- CP-element group 356: 	210 
    -- CP-element group 356:  members (15) 
      -- CP-element group 356: 	 branch_block_stmt_1049/if_stmt_2033__entry__
      -- CP-element group 356: 	 branch_block_stmt_1049/merge_stmt_2012__exit__
      -- CP-element group 356: 	 branch_block_stmt_1049/assign_stmt_2026_to_assign_stmt_2032__entry__
      -- CP-element group 356: 	 branch_block_stmt_1049/assign_stmt_2026_to_assign_stmt_2032__exit__
      -- CP-element group 356: 	 branch_block_stmt_1049/assign_stmt_2026_to_assign_stmt_2032/$entry
      -- CP-element group 356: 	 branch_block_stmt_1049/assign_stmt_2026_to_assign_stmt_2032/$exit
      -- CP-element group 356: 	 branch_block_stmt_1049/if_stmt_2033_dead_link/$entry
      -- CP-element group 356: 	 branch_block_stmt_1049/if_stmt_2033_eval_test/$entry
      -- CP-element group 356: 	 branch_block_stmt_1049/if_stmt_2033_eval_test/$exit
      -- CP-element group 356: 	 branch_block_stmt_1049/if_stmt_2033_eval_test/branch_req
      -- CP-element group 356: 	 branch_block_stmt_1049/R_tobool218_2034_place
      -- CP-element group 356: 	 branch_block_stmt_1049/if_stmt_2033_if_link/$entry
      -- CP-element group 356: 	 branch_block_stmt_1049/if_stmt_2033_else_link/$entry
      -- CP-element group 356: 	 branch_block_stmt_1049/merge_stmt_2012_PhiAck/$exit
      -- CP-element group 356: 	 branch_block_stmt_1049/merge_stmt_2012_PhiAck/phi_stmt_2013_ack
      -- 
    phi_stmt_2013_ack_6005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2013_ack_0, ack => convolution3D_CP_3189_elements(356)); -- 
    branch_req_4897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(356), ack => if_stmt_2033_branch_req_0); -- 
    -- CP-element group 357:  transition  output  delay-element  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	212 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (4) 
      -- CP-element group 357: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/$exit
      -- CP-element group 357: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/$exit
      -- CP-element group 357: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2071_konst_delay_trans
      -- CP-element group 357: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_req
      -- 
    phi_stmt_2065_req_6028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2065_req_6028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(357), ack => phi_stmt_2065_req_1); -- 
    -- Element group convolution3D_CP_3189_elements(357) is a control-delay.
    cp_element_357_delay: control_delay_element  generic map(name => " 357_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(212), ack => convolution3D_CP_3189_elements(357), clk => clk, reset =>reset);
    -- CP-element group 358:  transition  output  delay-element  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	212 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (4) 
      -- CP-element group 358: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/$exit
      -- CP-element group 358: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$exit
      -- CP-element group 358: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2064_konst_delay_trans
      -- CP-element group 358: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_req
      -- 
    phi_stmt_2058_req_6036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2058_req_6036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(358), ack => phi_stmt_2058_req_1); -- 
    -- Element group convolution3D_CP_3189_elements(358) is a control-delay.
    cp_element_358_delay: control_delay_element  generic map(name => " 358_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(212), ack => convolution3D_CP_3189_elements(358), clk => clk, reset =>reset);
    -- CP-element group 359:  join  transition  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	367 
    -- CP-element group 359:  members (1) 
      -- CP-element group 359: 	 branch_block_stmt_1049/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(357) & convolution3D_CP_3189_elements(358);
      gj_convolution3D_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	220 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (2) 
      -- CP-element group 360: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Sample/ra
      -- 
    ra_6056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2068_inst_ack_0, ack => convolution3D_CP_3189_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	220 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (2) 
      -- CP-element group 361: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/Update/ca
      -- 
    ca_6061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2068_inst_ack_1, ack => convolution3D_CP_3189_elements(361)); -- 
    -- CP-element group 362:  join  transition  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	366 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/$exit
      -- CP-element group 362: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/$exit
      -- CP-element group 362: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/$exit
      -- CP-element group 362: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_sources/type_cast_2068/SplitProtocol/$exit
      -- CP-element group 362: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2065/phi_stmt_2065_req
      -- 
    phi_stmt_2065_req_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2065_req_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(362), ack => phi_stmt_2065_req_0); -- 
    convolution3D_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(360) & convolution3D_CP_3189_elements(361);
      gj_convolution3D_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	220 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (2) 
      -- CP-element group 363: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/ra
      -- 
    ra_6079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_0, ack => convolution3D_CP_3189_elements(363)); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	220 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (2) 
      -- CP-element group 364: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/ca
      -- 
    ca_6084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_1, ack => convolution3D_CP_3189_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (5) 
      -- CP-element group 365: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/$exit
      -- CP-element group 365: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$exit
      -- CP-element group 365: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/$exit
      -- CP-element group 365: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/$exit
      -- CP-element group 365: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2058/phi_stmt_2058_req
      -- 
    phi_stmt_2058_req_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2058_req_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(365), ack => phi_stmt_2058_req_0); -- 
    convolution3D_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(363) & convolution3D_CP_3189_elements(364);
      gj_convolution3D_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	362 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (1) 
      -- CP-element group 366: 	 branch_block_stmt_1049/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(362) & convolution3D_CP_3189_elements(365);
      gj_convolution3D_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  merge  fork  transition  place  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	359 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_1049/merge_stmt_2057_PhiReqMerge
      -- CP-element group 367: 	 branch_block_stmt_1049/merge_stmt_2057_PhiAck/$entry
      -- 
    convolution3D_CP_3189_elements(367) <= OrReduce(convolution3D_CP_3189_elements(359) & convolution3D_CP_3189_elements(366));
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (1) 
      -- CP-element group 368: 	 branch_block_stmt_1049/merge_stmt_2057_PhiAck/phi_stmt_2058_ack
      -- 
    phi_stmt_2058_ack_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2058_ack_0, ack => convolution3D_CP_3189_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (1) 
      -- CP-element group 369: 	 branch_block_stmt_1049/merge_stmt_2057_PhiAck/phi_stmt_2065_ack
      -- 
    phi_stmt_2065_ack_6091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2065_ack_0, ack => convolution3D_CP_3189_elements(369)); -- 
    -- CP-element group 370:  join  fork  transition  place  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	213 
    -- CP-element group 370: 	216 
    -- CP-element group 370: 	217 
    -- CP-element group 370: 	218 
    -- CP-element group 370:  members (16) 
      -- CP-element group 370: 	 branch_block_stmt_1049/merge_stmt_2057__exit__
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111__entry__
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/$entry
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/RPIPE_maxpool_input_pipe_2086_Sample/rr
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_update_start_
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2090_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_update_start_
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Sample/rr
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_1049/assign_stmt_2078_to_assign_stmt_2111/type_cast_2105_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_1049/merge_stmt_2057_PhiAck/$exit
      -- 
    rr_4936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(370), ack => RPIPE_maxpool_input_pipe_2086_inst_req_0); -- 
    cr_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(370), ack => type_cast_2090_inst_req_1); -- 
    rr_4964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(370), ack => type_cast_2105_inst_req_0); -- 
    cr_4969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(370), ack => type_cast_2105_inst_req_1); -- 
    convolution3D_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(368) & convolution3D_CP_3189_elements(369);
      gj_convolution3D_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	221 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Sample/ra
      -- 
    ra_6115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2122_inst_ack_0, ack => convolution3D_CP_3189_elements(371)); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	221 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (2) 
      -- CP-element group 372: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/Update/ca
      -- 
    ca_6120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2122_inst_ack_1, ack => convolution3D_CP_3189_elements(372)); -- 
    -- CP-element group 373:  join  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (8) 
      -- CP-element group 373: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$exit
      -- CP-element group 373: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/$exit
      -- CP-element group 373: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/$exit
      -- CP-element group 373: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/$exit
      -- CP-element group 373: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_sources/type_cast_2122/SplitProtocol/$exit
      -- CP-element group 373: 	 branch_block_stmt_1049/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2119/phi_stmt_2119_req
      -- CP-element group 373: 	 branch_block_stmt_1049/merge_stmt_2118_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_1049/merge_stmt_2118_PhiAck/$entry
      -- 
    phi_stmt_2119_req_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2119_req_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(373), ack => phi_stmt_2119_req_0); -- 
    convolution3D_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(371) & convolution3D_CP_3189_elements(372);
      gj_convolution3D_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	227 
    -- CP-element group 374: 	222 
    -- CP-element group 374: 	223 
    -- CP-element group 374: 	225 
    -- CP-element group 374:  members (29) 
      -- CP-element group 374: 	 branch_block_stmt_1049/merge_stmt_2118__exit__
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157__entry__
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_update_start_
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_resized_1
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_scaled_1
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_computed_1
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_resize_1/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_resize_1/$exit
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_resize_1/index_resize_req
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_resize_1/index_resize_ack
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_scale_1/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_scale_1/$exit
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_scale_1/scale_rename_req
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_index_scale_1/scale_rename_ack
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_update_start
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Sample/req
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/array_obj_ref_2151_final_index_sum_regn_Update/req
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_complete/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/addr_of_2152_complete/req
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_update_start_
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/word_access_complete/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/word_access_complete/word_0/$entry
      -- CP-element group 374: 	 branch_block_stmt_1049/assign_stmt_2129_to_assign_stmt_2157/ptr_deref_2155_Update/word_access_complete/word_0/cr
      -- CP-element group 374: 	 branch_block_stmt_1049/merge_stmt_2118_PhiAck/$exit
      -- CP-element group 374: 	 branch_block_stmt_1049/merge_stmt_2118_PhiAck/phi_stmt_2119_ack
      -- 
    phi_stmt_2119_ack_6126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2119_ack_0, ack => convolution3D_CP_3189_elements(374)); -- 
    req_5017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(374), ack => array_obj_ref_2151_index_offset_req_0); -- 
    req_5022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(374), ack => array_obj_ref_2151_index_offset_req_1); -- 
    req_5037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(374), ack => addr_of_2152_final_reg_req_1); -- 
    cr_5087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(374), ack => ptr_deref_2155_store_0_req_1); -- 
    -- CP-element group 375:  merge  place  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	228 
    -- CP-element group 375: 	209 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (1) 
      -- CP-element group 375: 	 branch_block_stmt_1049/merge_stmt_2159_PhiReqMerge
      -- 
    convolution3D_CP_3189_elements(375) <= OrReduce(convolution3D_CP_3189_elements(228) & convolution3D_CP_3189_elements(209));
    -- CP-element group 376:  join  fork  transition  place  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	229 
    -- CP-element group 376: 	230 
    -- CP-element group 376:  members (36) 
      -- CP-element group 376: 	 branch_block_stmt_1049/merge_stmt_2159__exit__
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172__entry__
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_update_start_
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_word_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_root_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_address_resized
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_addr_resize/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_addr_resize/$exit
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_addr_resize/base_resize_req
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_addr_resize/base_resize_ack
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_plus_offset/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_plus_offset/$exit
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_plus_offset/sum_rename_req
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_base_plus_offset/sum_rename_ack
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_word_addrgen/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_word_addrgen/$exit
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_word_addrgen/root_register_req
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_word_addrgen/root_register_ack
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/ptr_deref_2169_Split/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/ptr_deref_2169_Split/$exit
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/ptr_deref_2169_Split/split_req
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/ptr_deref_2169_Split/split_ack
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/word_access_start/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/word_access_start/word_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Sample/word_access_start/word_0/rr
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/word_access_complete/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/word_access_complete/word_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/assign_stmt_2167_to_assign_stmt_2172/ptr_deref_2169_Update/word_access_complete/word_0/cr
      -- CP-element group 376: 	 branch_block_stmt_1049/merge_stmt_2159_PhiAck/$entry
      -- CP-element group 376: 	 branch_block_stmt_1049/merge_stmt_2159_PhiAck/$exit
      -- CP-element group 376: 	 branch_block_stmt_1049/merge_stmt_2159_PhiAck/dummy
      -- 
    rr_5129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(376), ack => ptr_deref_2169_store_0_req_0); -- 
    cr_5140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(376), ack => ptr_deref_2169_store_0_req_1); -- 
    convolution3D_CP_3189_elements(376) <= convolution3D_CP_3189_elements(375);
    -- CP-element group 377:  transition  output  delay-element  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	244 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	381 
    -- CP-element group 377:  members (5) 
      -- CP-element group 377: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- CP-element group 377: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2218/$exit
      -- CP-element group 377: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/$exit
      -- CP-element group 377: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2222_konst_delay_trans
      -- CP-element group 377: 	 branch_block_stmt_1049/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_req
      -- 
    phi_stmt_2218_req_6148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2218_req_6148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(377), ack => phi_stmt_2218_req_0); -- 
    -- Element group convolution3D_CP_3189_elements(377) is a control-delay.
    cp_element_377_delay: control_delay_element  generic map(name => " 377_delay", delay_value => 1)  port map(req => convolution3D_CP_3189_elements(244), ack => convolution3D_CP_3189_elements(377), clk => clk, reset =>reset);
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	255 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Sample/ra
      -- 
    ra_6168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2224_inst_ack_0, ack => convolution3D_CP_3189_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	255 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (2) 
      -- CP-element group 379: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/Update/ca
      -- 
    ca_6173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2224_inst_ack_1, ack => convolution3D_CP_3189_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (6) 
      -- CP-element group 380: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 380: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/$exit
      -- CP-element group 380: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/$exit
      -- CP-element group 380: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/$exit
      -- CP-element group 380: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2224/SplitProtocol/$exit
      -- CP-element group 380: 	 branch_block_stmt_1049/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2218/phi_stmt_2218_req
      -- 
    phi_stmt_2218_req_6174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2218_req_6174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(380), ack => phi_stmt_2218_req_1); -- 
    convolution3D_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3189_elements(378) & convolution3D_CP_3189_elements(379);
      gj_convolution3D_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3189_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  merge  transition  place  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	377 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (2) 
      -- CP-element group 381: 	 branch_block_stmt_1049/merge_stmt_2217_PhiReqMerge
      -- CP-element group 381: 	 branch_block_stmt_1049/merge_stmt_2217_PhiAck/$entry
      -- 
    convolution3D_CP_3189_elements(381) <= OrReduce(convolution3D_CP_3189_elements(377) & convolution3D_CP_3189_elements(380));
    -- CP-element group 382:  fork  transition  place  input  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	249 
    -- CP-element group 382: 	250 
    -- CP-element group 382: 	251 
    -- CP-element group 382: 	252 
    -- CP-element group 382: 	245 
    -- CP-element group 382:  members (20) 
      -- CP-element group 382: 	 branch_block_stmt_1049/merge_stmt_2217__exit__
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260__entry__
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_sample_start_
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_update_start_
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Sample/crr
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Sample/req
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/WPIPE_num_out_pipe_2231_sample_start_
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/$entry
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Update/ccr
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Sample/crr
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_update_start_
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2249_sample_start_
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_1049/assign_stmt_2230_to_assign_stmt_2260/call_stmt_2245_Update/ccr
      -- CP-element group 382: 	 branch_block_stmt_1049/merge_stmt_2217_PhiAck/$exit
      -- CP-element group 382: 	 branch_block_stmt_1049/merge_stmt_2217_PhiAck/phi_stmt_2218_ack
      -- 
    phi_stmt_2218_ack_6179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2218_ack_0, ack => convolution3D_CP_3189_elements(382)); -- 
    crr_5270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(382), ack => call_stmt_2245_call_req_0); -- 
    req_5242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(382), ack => WPIPE_num_out_pipe_2231_inst_req_0); -- 
    ccr_5289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(382), ack => call_stmt_2249_call_req_1); -- 
    crr_5284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(382), ack => call_stmt_2249_call_req_0); -- 
    ccr_5275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3189_elements(382), ack => call_stmt_2245_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1547_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1734_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_2008_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_2323_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1664 : std_logic_vector(63 downto 0);
    signal R_indvar411_1830_resized : std_logic_vector(13 downto 0);
    signal R_indvar411_1830_scaled : std_logic_vector(13 downto 0);
    signal R_indvar425_1369_resized : std_logic_vector(13 downto 0);
    signal R_indvar425_1369_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1685_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1685_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2150_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2150_scaled : std_logic_vector(13 downto 0);
    signal add102_1415 : std_logic_vector(63 downto 0);
    signal add108_1433 : std_logic_vector(63 downto 0);
    signal add114_1451 : std_logic_vector(63 downto 0);
    signal add120_1469 : std_logic_vector(63 downto 0);
    signal add1216x_xi370_2135 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1670 : std_logic_vector(63 downto 0);
    signal add126_1487 : std_logic_vector(63 downto 0);
    signal add132_1505 : std_logic_vector(63 downto 0);
    signal add13_1100 : std_logic_vector(15 downto 0);
    signal add171_1858 : std_logic_vector(63 downto 0);
    signal add177_1876 : std_logic_vector(63 downto 0);
    signal add183_1894 : std_logic_vector(63 downto 0);
    signal add189_1912 : std_logic_vector(63 downto 0);
    signal add195_1930 : std_logic_vector(63 downto 0);
    signal add201_1948 : std_logic_vector(63 downto 0);
    signal add207_1966 : std_logic_vector(63 downto 0);
    signal add23_1125 : std_logic_vector(15 downto 0);
    signal add33_1150 : std_logic_vector(15 downto 0);
    signal add43_1175 : std_logic_vector(15 downto 0);
    signal add53_1200 : std_logic_vector(15 downto 0);
    signal add63_1225 : std_logic_vector(63 downto 0);
    signal add73_1250 : std_logic_vector(15 downto 0);
    signal add96_1397 : std_logic_vector(63 downto 0);
    signal add_1075 : std_logic_vector(31 downto 0);
    signal addx_xi361_2096 : std_logic_vector(63 downto 0);
    signal addx_xi_1631 : std_logic_vector(63 downto 0);
    signal and217_2026 : std_logic_vector(63 downto 0);
    signal and_1565 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1370_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1370_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1370_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1370_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1370_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1370_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1831_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1831_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1831_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1831_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1831_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1831_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2151_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2151_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2151_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2151_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2151_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2151_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1688 : std_logic_vector(31 downto 0);
    signal arrayidx211_1833 : std_logic_vector(31 downto 0);
    signal arrayidx226_2153 : std_logic_vector(31 downto 0);
    signal arrayidx_1372 : std_logic_vector(31 downto 0);
    signal call105_1424 : std_logic_vector(7 downto 0);
    signal call111_1442 : std_logic_vector(7 downto 0);
    signal call117_1460 : std_logic_vector(7 downto 0);
    signal call11_1091 : std_logic_vector(7 downto 0);
    signal call123_1478 : std_logic_vector(7 downto 0);
    signal call129_1496 : std_logic_vector(7 downto 0);
    signal call164_1836 : std_logic_vector(7 downto 0);
    signal call168_1849 : std_logic_vector(7 downto 0);
    signal call16_1103 : std_logic_vector(7 downto 0);
    signal call174_1867 : std_logic_vector(7 downto 0);
    signal call180_1885 : std_logic_vector(7 downto 0);
    signal call186_1903 : std_logic_vector(7 downto 0);
    signal call192_1921 : std_logic_vector(7 downto 0);
    signal call198_1939 : std_logic_vector(7 downto 0);
    signal call204_1957 : std_logic_vector(7 downto 0);
    signal call21_1116 : std_logic_vector(7 downto 0);
    signal call229_2175 : std_logic_vector(63 downto 0);
    signal call26_1128 : std_logic_vector(7 downto 0);
    signal call270_2275 : std_logic_vector(7 downto 0);
    signal call273_2279 : std_logic_vector(7 downto 0);
    signal call275_2282 : std_logic_vector(63 downto 0);
    signal call2_1066 : std_logic_vector(7 downto 0);
    signal call31_1141 : std_logic_vector(7 downto 0);
    signal call36_1153 : std_logic_vector(7 downto 0);
    signal call41_1166 : std_logic_vector(7 downto 0);
    signal call46_1178 : std_logic_vector(7 downto 0);
    signal call51_1191 : std_logic_vector(7 downto 0);
    signal call56_1203 : std_logic_vector(7 downto 0);
    signal call61_1216 : std_logic_vector(7 downto 0);
    signal call66_1228 : std_logic_vector(7 downto 0);
    signal call6_1078 : std_logic_vector(7 downto 0);
    signal call71_1241 : std_logic_vector(7 downto 0);
    signal call89_1375 : std_logic_vector(7 downto 0);
    signal call93_1388 : std_logic_vector(7 downto 0);
    signal call99_1406 : std_logic_vector(7 downto 0);
    signal call_1053 : std_logic_vector(7 downto 0);
    signal callx_xi359_2087 : std_logic_vector(7 downto 0);
    signal callx_xi_1622 : std_logic_vector(7 downto 0);
    signal cmp161379_1742 : std_logic_vector(0 downto 0);
    signal cmp383_1279 : std_logic_vector(0 downto 0);
    signal cmpx_xi364_2111 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1646 : std_logic_vector(0 downto 0);
    signal conv101_1410 : std_logic_vector(63 downto 0);
    signal conv107_1428 : std_logic_vector(63 downto 0);
    signal conv113_1446 : std_logic_vector(63 downto 0);
    signal conv119_1464 : std_logic_vector(63 downto 0);
    signal conv125_1482 : std_logic_vector(63 downto 0);
    signal conv12_1095 : std_logic_vector(15 downto 0);
    signal conv131_1500 : std_logic_vector(63 downto 0);
    signal conv145_1698 : std_logic_vector(63 downto 0);
    signal conv147_1702 : std_logic_vector(63 downto 0);
    signal conv153_1706 : std_logic_vector(63 downto 0);
    signal conv155_1736 : std_logic_vector(63 downto 0);
    signal conv165_1840 : std_logic_vector(63 downto 0);
    signal conv170_1853 : std_logic_vector(63 downto 0);
    signal conv176_1871 : std_logic_vector(63 downto 0);
    signal conv182_1889 : std_logic_vector(63 downto 0);
    signal conv188_1907 : std_logic_vector(63 downto 0);
    signal conv194_1925 : std_logic_vector(63 downto 0);
    signal conv19_1107 : std_logic_vector(15 downto 0);
    signal conv1_1057 : std_logic_vector(31 downto 0);
    signal conv200_1943 : std_logic_vector(63 downto 0);
    signal conv206_1961 : std_logic_vector(63 downto 0);
    signal conv22_1120 : std_logic_vector(15 downto 0);
    signal conv230_2272 : std_logic_vector(63 downto 0);
    signal conv254_2242 : std_logic_vector(63 downto 0);
    signal conv276_2287 : std_logic_vector(63 downto 0);
    signal conv281_2296 : std_logic_vector(63 downto 0);
    signal conv283_2300 : std_logic_vector(63 downto 0);
    signal conv288_2325 : std_logic_vector(63 downto 0);
    signal conv292_2332 : std_logic_vector(7 downto 0);
    signal conv298_2342 : std_logic_vector(7 downto 0);
    signal conv29_1132 : std_logic_vector(15 downto 0);
    signal conv2x_xi354_2049 : std_logic_vector(31 downto 0);
    signal conv2x_xi_1584 : std_logic_vector(31 downto 0);
    signal conv304_2352 : std_logic_vector(7 downto 0);
    signal conv310_2362 : std_logic_vector(7 downto 0);
    signal conv316_2372 : std_logic_vector(7 downto 0);
    signal conv322_2382 : std_logic_vector(7 downto 0);
    signal conv328_2392 : std_logic_vector(7 downto 0);
    signal conv32_1145 : std_logic_vector(15 downto 0);
    signal conv334_2402 : std_logic_vector(7 downto 0);
    signal conv39_1157 : std_logic_vector(15 downto 0);
    signal conv3_1070 : std_logic_vector(31 downto 0);
    signal conv42_1170 : std_logic_vector(15 downto 0);
    signal conv49_1182 : std_logic_vector(15 downto 0);
    signal conv52_1195 : std_logic_vector(15 downto 0);
    signal conv59_1207 : std_logic_vector(63 downto 0);
    signal conv5x_xi360_2091 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1626 : std_logic_vector(63 downto 0);
    signal conv62_1220 : std_logic_vector(63 downto 0);
    signal conv69_1232 : std_logic_vector(15 downto 0);
    signal conv72_1245 : std_logic_vector(15 downto 0);
    signal conv79_1254 : std_logic_vector(31 downto 0);
    signal conv81_1258 : std_logic_vector(31 downto 0);
    signal conv83_1273 : std_logic_vector(63 downto 0);
    signal conv90_1379 : std_logic_vector(63 downto 0);
    signal conv95_1392 : std_logic_vector(63 downto 0);
    signal conv9_1082 : std_logic_vector(15 downto 0);
    signal convx_xi363_2106 : std_logic_vector(31 downto 0);
    signal convx_xi_1641 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi358_2065 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_1600 : std_logic_vector(63 downto 0);
    signal exitcond28_1520 : std_logic_vector(0 downto 0);
    signal exitcond5_2260 : std_logic_vector(0 downto 0);
    signal exitcond_1981 : std_logic_vector(0 downto 0);
    signal iNsTr_35_1619 : std_logic_vector(15 downto 0);
    signal iNsTr_48_2167 : std_logic_vector(31 downto 0);
    signal iNsTr_59_2045 : std_logic_vector(63 downto 0);
    signal iNsTr_71_2084 : std_logic_vector(15 downto 0);
    signal iNsTr_97_2129 : std_logic_vector(63 downto 0);
    signal indvar411_1819 : std_logic_vector(63 downto 0);
    signal indvar425_1358 : std_logic_vector(63 downto 0);
    signal indvar_2218 : std_logic_vector(63 downto 0);
    signal indvarx_xnext412_1976 : std_logic_vector(63 downto 0);
    signal indvarx_xnext426_1515 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_2255 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_1552 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_2013 : std_logic_vector(63 downto 0);
    signal mul148_1711 : std_logic_vector(63 downto 0);
    signal mul151_1716 : std_logic_vector(63 downto 0);
    signal mul154_1721 : std_logic_vector(63 downto 0);
    signal mul253_2230 : std_logic_vector(63 downto 0);
    signal mul284_2306 : std_logic_vector(63 downto 0);
    signal mul287_2311 : std_logic_vector(63 downto 0);
    signal mul82_1268 : std_logic_vector(31 downto 0);
    signal mul_1263 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi357_2058 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_1593 : std_logic_vector(15 downto 0);
    signal phitmp387_2010 : std_logic_vector(63 downto 0);
    signal phitmp_1549 : std_logic_vector(63 downto 0);
    signal ptr_deref_1507_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1507_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1507_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1507_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1507_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1507_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1690_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1690_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1690_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1690_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1690_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1690_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1968_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1968_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1968_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1968_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1968_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1968_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2155_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2155_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2155_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2155_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2155_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2155_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2169_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2169_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext352_2316 : std_logic_vector(63 downto 0);
    signal sext_1727 : std_logic_vector(63 downto 0);
    signal sh_promx_xi371_2141 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1676 : std_logic_vector(63 downto 0);
    signal shl104_1421 : std_logic_vector(63 downto 0);
    signal shl10_1088 : std_logic_vector(15 downto 0);
    signal shl110_1439 : std_logic_vector(63 downto 0);
    signal shl116_1457 : std_logic_vector(63 downto 0);
    signal shl122_1475 : std_logic_vector(63 downto 0);
    signal shl128_1493 : std_logic_vector(63 downto 0);
    signal shl14x_xi372_2146 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1681 : std_logic_vector(63 downto 0);
    signal shl167_1846 : std_logic_vector(63 downto 0);
    signal shl173_1864 : std_logic_vector(63 downto 0);
    signal shl179_1882 : std_logic_vector(63 downto 0);
    signal shl185_1900 : std_logic_vector(63 downto 0);
    signal shl191_1918 : std_logic_vector(63 downto 0);
    signal shl197_1936 : std_logic_vector(63 downto 0);
    signal shl203_1954 : std_logic_vector(63 downto 0);
    signal shl20_1113 : std_logic_vector(15 downto 0);
    signal shl30_1138 : std_logic_vector(15 downto 0);
    signal shl40_1163 : std_logic_vector(15 downto 0);
    signal shl50_1188 : std_logic_vector(15 downto 0);
    signal shl60_1213 : std_logic_vector(63 downto 0);
    signal shl70_1238 : std_logic_vector(15 downto 0);
    signal shl8x_xi362_2102 : std_logic_vector(63 downto 0);
    signal shl8x_xi362x_xlcssa_2119 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1637 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1654 : std_logic_vector(63 downto 0);
    signal shl92_1385 : std_logic_vector(63 downto 0);
    signal shl98_1403 : std_logic_vector(63 downto 0);
    signal shl_1063 : std_logic_vector(31 downto 0);
    signal shlx_xi355_2055 : std_logic_vector(31 downto 0);
    signal shlx_xi_1590 : std_logic_vector(31 downto 0);
    signal shr295_2338 : std_logic_vector(63 downto 0);
    signal shr301_2348 : std_logic_vector(63 downto 0);
    signal shr307_2358 : std_logic_vector(63 downto 0);
    signal shr313_2368 : std_logic_vector(63 downto 0);
    signal shr319_2378 : std_logic_vector(63 downto 0);
    signal shr325_2388 : std_logic_vector(63 downto 0);
    signal shr331_2398 : std_logic_vector(63 downto 0);
    signal sub_2292 : std_logic_vector(63 downto 0);
    signal tmp10_1770 : std_logic_vector(63 downto 0);
    signal tmp11_1774 : std_logic_vector(63 downto 0);
    signal tmp12_1779 : std_logic_vector(63 downto 0);
    signal tmp13_1783 : std_logic_vector(63 downto 0);
    signal tmp14_1788 : std_logic_vector(63 downto 0);
    signal tmp15_1792 : std_logic_vector(31 downto 0);
    signal tmp16_1797 : std_logic_vector(63 downto 0);
    signal tmp17_1803 : std_logic_vector(63 downto 0);
    signal tmp18_1809 : std_logic_vector(0 downto 0);
    signal tmp20_1317 : std_logic_vector(31 downto 0);
    signal tmp21_1322 : std_logic_vector(31 downto 0);
    signal tmp22_1326 : std_logic_vector(31 downto 0);
    signal tmp23_1331 : std_logic_vector(31 downto 0);
    signal tmp24_1336 : std_logic_vector(63 downto 0);
    signal tmp25_1342 : std_logic_vector(63 downto 0);
    signal tmp26_1348 : std_logic_vector(0 downto 0);
    signal tmp388_2078 : std_logic_vector(15 downto 0);
    signal tmp389_2191 : std_logic_vector(15 downto 0);
    signal tmp393_2196 : std_logic_vector(15 downto 0);
    signal tmp3_2200 : std_logic_vector(63 downto 0);
    signal tmp406_1755 : std_logic_vector(63 downto 0);
    signal tmp407_1761 : std_logic_vector(0 downto 0);
    signal tmp408_2001 : std_logic_vector(63 downto 0);
    signal tmp415_1291 : std_logic_vector(31 downto 0);
    signal tmp417_1296 : std_logic_vector(31 downto 0);
    signal tmp418_1301 : std_logic_vector(63 downto 0);
    signal tmp419_1307 : std_logic_vector(63 downto 0);
    signal tmp420_1313 : std_logic_vector(0 downto 0);
    signal tmp422_1540 : std_logic_vector(63 downto 0);
    signal tmp4_2206 : std_logic_vector(63 downto 0);
    signal tmp6_2210 : std_logic_vector(63 downto 0);
    signal tmp7_2215 : std_logic_vector(63 downto 0);
    signal tmp9_1765 : std_logic_vector(63 downto 0);
    signal tmp_1613 : std_logic_vector(15 downto 0);
    signal tobool218_2032 : std_logic_vector(0 downto 0);
    signal tobool_1571 : std_logic_vector(0 downto 0);
    signal type_cast_1061_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1086_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1111_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1136_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1161_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1186_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1211_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1271_wire : std_logic_vector(63 downto 0);
    signal type_cast_1277_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1299_wire : std_logic_vector(63 downto 0);
    signal type_cast_1305_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1311_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1334_wire : std_logic_vector(63 downto 0);
    signal type_cast_1340_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1346_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1353_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1362_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1364_wire : std_logic_vector(63 downto 0);
    signal type_cast_1383_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1401_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1419_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1437_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1455_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1473_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1491_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1538_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1543_wire : std_logic_vector(63 downto 0);
    signal type_cast_1546_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1555_wire : std_logic_vector(63 downto 0);
    signal type_cast_1558_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1563_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1569_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1582_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1588_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1597_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1599_wire : std_logic_vector(15 downto 0);
    signal type_cast_1604_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1606_wire : std_logic_vector(63 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1617_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1635_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1657_wire : std_logic_vector(63 downto 0);
    signal type_cast_1662_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1668_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1674_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1725_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1730_wire : std_logic_vector(63 downto 0);
    signal type_cast_1733_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1740_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1753_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1759_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1795_wire : std_logic_vector(63 downto 0);
    signal type_cast_1801_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1807_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1814_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1822_wire : std_logic_vector(63 downto 0);
    signal type_cast_1825_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1844_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1862_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1880_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1898_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1916_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1934_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1952_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1974_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1993_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1999_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2004_wire : std_logic_vector(63 downto 0);
    signal type_cast_2007_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2016_wire : std_logic_vector(63 downto 0);
    signal type_cast_2019_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2024_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2043_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2053_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2061_wire : std_logic_vector(15 downto 0);
    signal type_cast_2064_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2068_wire : std_logic_vector(63 downto 0);
    signal type_cast_2071_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2076_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2082_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2100_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2122_wire : std_logic_vector(63 downto 0);
    signal type_cast_2127_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2133_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2139_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2171_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2189_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2204_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2222_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2224_wire : std_logic_vector(63 downto 0);
    signal type_cast_2240_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2253_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2270_wire : std_logic_vector(63 downto 0);
    signal type_cast_2285_wire : std_logic_vector(63 downto 0);
    signal type_cast_2304_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2319_wire : std_logic_vector(63 downto 0);
    signal type_cast_2322_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2336_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2346_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2356_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2366_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2376_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2386_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2396_wire_constant : std_logic_vector(63 downto 0);
    signal umax19_1816 : std_logic_vector(63 downto 0);
    signal umax27_1355 : std_logic_vector(63 downto 0);
    signal umax421_1534 : std_logic_vector(63 downto 0);
    signal umax_1995 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1370_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1370_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1370_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1370_resized_base_address <= "00000000000000";
    array_obj_ref_1686_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1686_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1686_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1686_resized_base_address <= "00000000000000";
    array_obj_ref_1831_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1831_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1831_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1831_resized_base_address <= "00000000000000";
    array_obj_ref_2151_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2151_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2151_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2151_resized_base_address <= "00000000000000";
    iNsTr_48_2167 <= "00000000000000000000000000000000";
    ptr_deref_1507_word_offset_0 <= "00000000000000";
    ptr_deref_1690_word_offset_0 <= "00000000000000";
    ptr_deref_1968_word_offset_0 <= "00000000000000";
    ptr_deref_2155_word_offset_0 <= "00000000000000";
    ptr_deref_2169_word_offset_0 <= "00000000000000";
    type_cast_1061_wire_constant <= "00000000000000000000000000001000";
    type_cast_1086_wire_constant <= "0000000000001000";
    type_cast_1111_wire_constant <= "0000000000001000";
    type_cast_1136_wire_constant <= "0000000000001000";
    type_cast_1161_wire_constant <= "0000000000001000";
    type_cast_1186_wire_constant <= "0000000000001000";
    type_cast_1211_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1236_wire_constant <= "0000000000001000";
    type_cast_1277_wire_constant <= "00000000000000000000000000000011";
    type_cast_1305_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1311_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1340_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1346_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1353_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1362_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1383_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1401_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1419_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1437_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1455_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1473_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1491_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1532_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1538_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1546_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1558_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1563_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1569_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1582_wire_constant <= "00000000000000000000000000000001";
    type_cast_1588_wire_constant <= "00000000000000000000000000000110";
    type_cast_1597_wire_constant <= "0000000000000000";
    type_cast_1604_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1611_wire_constant <= "0000000000000001";
    type_cast_1617_wire_constant <= "0000000000000001";
    type_cast_1635_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1662_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1668_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1674_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1725_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1733_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1740_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1753_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1759_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1801_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1807_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1814_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1825_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1844_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1862_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1880_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1898_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1916_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1934_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1952_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1974_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1993_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1999_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2007_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2019_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2024_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2043_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2053_wire_constant <= "00000000000000000000000000000110";
    type_cast_2064_wire_constant <= "0000000000000000";
    type_cast_2071_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2076_wire_constant <= "0000000000000001";
    type_cast_2082_wire_constant <= "0000000000000001";
    type_cast_2100_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2127_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_2133_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2139_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2171_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2189_wire_constant <= "1111111111111111";
    type_cast_2204_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2240_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_2253_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2304_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2322_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2336_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2346_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2356_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2366_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2376_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_1358: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1362_wire_constant & type_cast_1364_wire;
      req <= phi_stmt_1358_req_0 & phi_stmt_1358_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1358",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1358_ack_0,
          idata => idata,
          odata => indvar425_1358,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1358
    phi_stmt_1552: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1555_wire & type_cast_1558_wire_constant;
      req <= phi_stmt_1552_req_0 & phi_stmt_1552_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1552",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1552_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1552,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1552
    phi_stmt_1593: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1597_wire_constant & type_cast_1599_wire;
      req <= phi_stmt_1593_req_0 & phi_stmt_1593_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1593",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1593_ack_0,
          idata => idata,
          odata => nx_x022x_xi_1593,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1593
    phi_stmt_1600: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1604_wire_constant & type_cast_1606_wire;
      req <= phi_stmt_1600_req_0 & phi_stmt_1600_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1600",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1600_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_1600,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1600
    phi_stmt_1654: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1657_wire;
      req(0) <= phi_stmt_1654_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1654",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1654_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1654,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1654
    phi_stmt_1819: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1822_wire & type_cast_1825_wire_constant;
      req <= phi_stmt_1819_req_0 & phi_stmt_1819_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1819",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1819_ack_0,
          idata => idata,
          odata => indvar411_1819,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1819
    phi_stmt_2013: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2016_wire & type_cast_2019_wire_constant;
      req <= phi_stmt_2013_req_0 & phi_stmt_2013_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2013",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2013_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_2013,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2013
    phi_stmt_2058: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2061_wire & type_cast_2064_wire_constant;
      req <= phi_stmt_2058_req_0 & phi_stmt_2058_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2058",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2058_ack_0,
          idata => idata,
          odata => nx_x022x_xi357_2058,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2058
    phi_stmt_2065: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2068_wire & type_cast_2071_wire_constant;
      req <= phi_stmt_2065_req_0 & phi_stmt_2065_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2065",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2065_ack_0,
          idata => idata,
          odata => elementx_x021x_xi358_2065,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2065
    phi_stmt_2119: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2122_wire;
      req(0) <= phi_stmt_2119_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2119",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2119_ack_0,
          idata => idata,
          odata => shl8x_xi362x_xlcssa_2119,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2119
    phi_stmt_2218: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2222_wire_constant & type_cast_2224_wire;
      req <= phi_stmt_2218_req_0 & phi_stmt_2218_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2218",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2218_ack_0,
          idata => idata,
          odata => indvar_2218,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2218
    -- flow-through select operator MUX_1354_inst
    umax27_1355 <= tmp25_1342 when (tmp26_1348(0) /=  '0') else type_cast_1353_wire_constant;
    -- flow-through select operator MUX_1533_inst
    umax421_1534 <= tmp419_1307 when (tmp420_1313(0) /=  '0') else type_cast_1532_wire_constant;
    -- flow-through select operator MUX_1815_inst
    umax19_1816 <= tmp17_1803 when (tmp18_1809(0) /=  '0') else type_cast_1814_wire_constant;
    -- flow-through select operator MUX_1994_inst
    umax_1995 <= tmp406_1755 when (tmp407_1761(0) /=  '0') else type_cast_1993_wire_constant;
    addr_of_1371_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1371_final_reg_req_0;
      addr_of_1371_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1371_final_reg_req_1;
      addr_of_1371_final_reg_ack_1<= rack(0);
      addr_of_1371_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1371_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1370_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1687_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1687_final_reg_req_0;
      addr_of_1687_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1687_final_reg_req_1;
      addr_of_1687_final_reg_ack_1<= rack(0);
      addr_of_1687_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1687_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1686_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1832_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1832_final_reg_req_0;
      addr_of_1832_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1832_final_reg_req_1;
      addr_of_1832_final_reg_ack_1<= rack(0);
      addr_of_1832_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1832_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1831_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2152_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2152_final_reg_req_0;
      addr_of_2152_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2152_final_reg_req_1;
      addr_of_2152_final_reg_ack_1<= rack(0);
      addr_of_2152_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2152_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2151_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_2153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1056_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1056_inst_req_0;
      type_cast_1056_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1056_inst_req_1;
      type_cast_1056_inst_ack_1<= rack(0);
      type_cast_1056_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1056_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1053,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1069_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1069_inst_req_0;
      type_cast_1069_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1069_inst_req_1;
      type_cast_1069_inst_ack_1<= rack(0);
      type_cast_1069_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1069_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1070,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1081_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1081_inst_req_0;
      type_cast_1081_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1081_inst_req_1;
      type_cast_1081_inst_ack_1<= rack(0);
      type_cast_1081_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1081_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1078,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_1082,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1094_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1094_inst_req_0;
      type_cast_1094_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1094_inst_req_1;
      type_cast_1094_inst_ack_1<= rack(0);
      type_cast_1094_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1094_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_1091,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1106_inst_req_0;
      type_cast_1106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1106_inst_req_1;
      type_cast_1106_inst_ack_1<= rack(0);
      type_cast_1106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1119_inst_req_0;
      type_cast_1119_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1119_inst_req_1;
      type_cast_1119_inst_ack_1<= rack(0);
      type_cast_1119_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_1116,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1131_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1131_inst_req_0;
      type_cast_1131_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1131_inst_req_1;
      type_cast_1131_inst_ack_1<= rack(0);
      type_cast_1131_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1131_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1144_inst_req_0;
      type_cast_1144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1144_inst_req_1;
      type_cast_1144_inst_ack_1<= rack(0);
      type_cast_1144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_1141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1156_inst_req_0;
      type_cast_1156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1156_inst_req_1;
      type_cast_1156_inst_ack_1<= rack(0);
      type_cast_1156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1169_inst_req_0;
      type_cast_1169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1169_inst_req_1;
      type_cast_1169_inst_ack_1<= rack(0);
      type_cast_1169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_1166,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1181_inst_req_0;
      type_cast_1181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1181_inst_req_1;
      type_cast_1181_inst_ack_1<= rack(0);
      type_cast_1181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_1178,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1194_inst_req_0;
      type_cast_1194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1194_inst_req_1;
      type_cast_1194_inst_ack_1<= rack(0);
      type_cast_1194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_1191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1206_inst_req_0;
      type_cast_1206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1206_inst_req_1;
      type_cast_1206_inst_ack_1<= rack(0);
      type_cast_1206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_1203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1219_inst_req_0;
      type_cast_1219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1219_inst_req_1;
      type_cast_1219_inst_ack_1<= rack(0);
      type_cast_1219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_1216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1231_inst_req_0;
      type_cast_1231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1231_inst_req_1;
      type_cast_1231_inst_ack_1<= rack(0);
      type_cast_1231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_1228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1244_inst_req_0;
      type_cast_1244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1244_inst_req_1;
      type_cast_1244_inst_ack_1<= rack(0);
      type_cast_1244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_1241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_1245,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1253_inst_req_0;
      type_cast_1253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1253_inst_req_1;
      type_cast_1253_inst_ack_1<= rack(0);
      type_cast_1253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1257_inst_req_0;
      type_cast_1257_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1257_inst_req_1;
      type_cast_1257_inst_ack_1<= rack(0);
      type_cast_1257_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1257_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1272_inst_req_0;
      type_cast_1272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1272_inst_req_1;
      type_cast_1272_inst_ack_1<= rack(0);
      type_cast_1272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1271_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1273,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1300_inst_req_0;
      type_cast_1300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1300_inst_req_1;
      type_cast_1300_inst_ack_1<= rack(0);
      type_cast_1300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1300_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1299_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp418_1301,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1316_inst_req_0;
      type_cast_1316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1316_inst_req_1;
      type_cast_1316_inst_ack_1<= rack(0);
      type_cast_1316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1325_inst_req_0;
      type_cast_1325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1325_inst_req_1;
      type_cast_1325_inst_ack_1<= rack(0);
      type_cast_1325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp22_1326,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1335_inst_req_0;
      type_cast_1335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1335_inst_req_1;
      type_cast_1335_inst_ack_1<= rack(0);
      type_cast_1335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1334_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_1336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1364_inst_req_0;
      type_cast_1364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1364_inst_req_1;
      type_cast_1364_inst_ack_1<= rack(0);
      type_cast_1364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext426_1515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1364_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1378_inst_req_0;
      type_cast_1378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1378_inst_req_1;
      type_cast_1378_inst_ack_1<= rack(0);
      type_cast_1378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_1375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1391_inst_req_0;
      type_cast_1391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1391_inst_req_1;
      type_cast_1391_inst_ack_1<= rack(0);
      type_cast_1391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_1388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_1392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1409_inst_req_0;
      type_cast_1409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1409_inst_req_1;
      type_cast_1409_inst_ack_1<= rack(0);
      type_cast_1409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_1406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_1410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1427_inst_req_0;
      type_cast_1427_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1427_inst_req_1;
      type_cast_1427_inst_ack_1<= rack(0);
      type_cast_1427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_1424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1445_inst_req_0;
      type_cast_1445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1445_inst_req_1;
      type_cast_1445_inst_ack_1<= rack(0);
      type_cast_1445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_1442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_1446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1463_inst_req_0;
      type_cast_1463_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1463_inst_req_1;
      type_cast_1463_inst_ack_1<= rack(0);
      type_cast_1463_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1463_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_1460,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_1464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1481_inst_req_0;
      type_cast_1481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1481_inst_req_1;
      type_cast_1481_inst_ack_1<= rack(0);
      type_cast_1481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_1478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_1482,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1499_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1499_inst_req_0;
      type_cast_1499_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1499_inst_req_1;
      type_cast_1499_inst_ack_1<= rack(0);
      type_cast_1499_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1499_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_1496,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_1500,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1543_inst
    process(tmp422_1540) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp422_1540(63 downto 0);
      type_cast_1543_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1548_inst
    process(ASHR_i64_i64_1547_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1547_wire(63 downto 0);
      phitmp_1549 <= tmp_var; -- 
    end process;
    type_cast_1555_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1555_inst_req_0;
      type_cast_1555_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1555_inst_req_1;
      type_cast_1555_inst_ack_1<= rack(0);
      type_cast_1555_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1555_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_1549,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1555_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1599_inst_req_0;
      type_cast_1599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1599_inst_req_1;
      type_cast_1599_inst_ack_1<= rack(0);
      type_cast_1599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_1619,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1599_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1606_inst_req_0;
      type_cast_1606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1606_inst_req_1;
      type_cast_1606_inst_ack_1<= rack(0);
      type_cast_1606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1637,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1606_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1625_inst_req_0;
      type_cast_1625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1625_inst_req_1;
      type_cast_1625_inst_ack_1<= rack(0);
      type_cast_1625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1626,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1640_inst_req_0;
      type_cast_1640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1640_inst_req_1;
      type_cast_1640_inst_ack_1<= rack(0);
      type_cast_1640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1641,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1657_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1657_inst_req_0;
      type_cast_1657_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1657_inst_req_1;
      type_cast_1657_inst_ack_1<= rack(0);
      type_cast_1657_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1657_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1637,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1657_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1697_inst_req_0;
      type_cast_1697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1697_inst_req_1;
      type_cast_1697_inst_ack_1<= rack(0);
      type_cast_1697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1701_inst_req_0;
      type_cast_1701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1701_inst_req_1;
      type_cast_1701_inst_ack_1<= rack(0);
      type_cast_1701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1705_inst_req_0;
      type_cast_1705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1705_inst_req_1;
      type_cast_1705_inst_ack_1<= rack(0);
      type_cast_1705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1730_inst
    process(sext_1727) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1727(63 downto 0);
      type_cast_1730_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1735_inst
    process(ASHR_i64_i64_1734_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1734_wire(63 downto 0);
      conv155_1736 <= tmp_var; -- 
    end process;
    type_cast_1764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1764_inst_req_0;
      type_cast_1764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1764_inst_req_1;
      type_cast_1764_inst_ack_1<= rack(0);
      type_cast_1764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp9_1765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1773_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1773_inst_req_0;
      type_cast_1773_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1773_inst_req_1;
      type_cast_1773_inst_ack_1<= rack(0);
      type_cast_1773_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1773_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp11_1774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1782_inst_req_0;
      type_cast_1782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1782_inst_req_1;
      type_cast_1782_inst_ack_1<= rack(0);
      type_cast_1782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1791_inst_req_0;
      type_cast_1791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1791_inst_req_1;
      type_cast_1791_inst_ack_1<= rack(0);
      type_cast_1791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_1788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1792,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1796_inst_req_0;
      type_cast_1796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1796_inst_req_1;
      type_cast_1796_inst_ack_1<= rack(0);
      type_cast_1796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1796_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1795_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_1797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1822_inst_req_0;
      type_cast_1822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1822_inst_req_1;
      type_cast_1822_inst_ack_1<= rack(0);
      type_cast_1822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext412_1976,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1822_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1839_inst_req_0;
      type_cast_1839_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1839_inst_req_1;
      type_cast_1839_inst_ack_1<= rack(0);
      type_cast_1839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1836,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1852_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1852_inst_req_0;
      type_cast_1852_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1852_inst_req_1;
      type_cast_1852_inst_ack_1<= rack(0);
      type_cast_1852_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1852_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1849,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1853,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1870_inst_req_0;
      type_cast_1870_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1870_inst_req_1;
      type_cast_1870_inst_ack_1<= rack(0);
      type_cast_1870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1867,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1871,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1888_inst_req_0;
      type_cast_1888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1888_inst_req_1;
      type_cast_1888_inst_ack_1<= rack(0);
      type_cast_1888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1888_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1885,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1889,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1906_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1906_inst_req_0;
      type_cast_1906_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1906_inst_req_1;
      type_cast_1906_inst_ack_1<= rack(0);
      type_cast_1906_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1906_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1903,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1907,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1924_inst_req_0;
      type_cast_1924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1924_inst_req_1;
      type_cast_1924_inst_ack_1<= rack(0);
      type_cast_1924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1921,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1942_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1942_inst_req_0;
      type_cast_1942_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1942_inst_req_1;
      type_cast_1942_inst_ack_1<= rack(0);
      type_cast_1942_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1942_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_1939,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_1943,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1960_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1960_inst_req_0;
      type_cast_1960_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1960_inst_req_1;
      type_cast_1960_inst_ack_1<= rack(0);
      type_cast_1960_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1960_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_1957,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_1961,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2004_inst
    process(tmp408_2001) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp408_2001(63 downto 0);
      type_cast_2004_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2009_inst
    process(ASHR_i64_i64_2008_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_2008_wire(63 downto 0);
      phitmp387_2010 <= tmp_var; -- 
    end process;
    type_cast_2016_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2016_inst_req_0;
      type_cast_2016_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2016_inst_req_1;
      type_cast_2016_inst_ack_1<= rack(0);
      type_cast_2016_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2016_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp387_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2016_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2048_inst_req_0;
      type_cast_2048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2048_inst_req_1;
      type_cast_2048_inst_ack_1<= rack(0);
      type_cast_2048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_59_2045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi354_2049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2061_inst_req_0;
      type_cast_2061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2061_inst_req_1;
      type_cast_2061_inst_ack_1<= rack(0);
      type_cast_2061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_71_2084,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2061_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2068_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2068_inst_req_0;
      type_cast_2068_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2068_inst_req_1;
      type_cast_2068_inst_ack_1<= rack(0);
      type_cast_2068_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2068_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_2102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2068_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2090_inst_req_0;
      type_cast_2090_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2090_inst_req_1;
      type_cast_2090_inst_ack_1<= rack(0);
      type_cast_2090_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2090_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi359_2087,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi360_2091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2105_inst_req_0;
      type_cast_2105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2105_inst_req_1;
      type_cast_2105_inst_ack_1<= rack(0);
      type_cast_2105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp388_2078,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi363_2106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2122_inst_req_0;
      type_cast_2122_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2122_inst_req_1;
      type_cast_2122_inst_ack_1<= rack(0);
      type_cast_2122_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2122_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_2102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2122_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2199_inst_req_0;
      type_cast_2199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2199_inst_req_1;
      type_cast_2199_inst_ack_1<= rack(0);
      type_cast_2199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp389_2191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_2200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2209_inst_req_0;
      type_cast_2209_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2209_inst_req_1;
      type_cast_2209_inst_ack_1<= rack(0);
      type_cast_2209_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2209_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp393_2196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_2210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2224_inst_req_0;
      type_cast_2224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2224_inst_req_1;
      type_cast_2224_inst_ack_1<= rack(0);
      type_cast_2224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2224_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2271_inst_req_0;
      type_cast_2271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2271_inst_req_1;
      type_cast_2271_inst_ack_1<= rack(0);
      type_cast_2271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2271_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2270_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_2272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2286_inst_req_0;
      type_cast_2286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2286_inst_req_1;
      type_cast_2286_inst_ack_1<= rack(0);
      type_cast_2286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2285_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_2287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2295_inst_req_0;
      type_cast_2295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2295_inst_req_1;
      type_cast_2295_inst_ack_1<= rack(0);
      type_cast_2295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add43_1175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv281_2296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2299_inst_req_0;
      type_cast_2299_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2299_inst_req_1;
      type_cast_2299_inst_ack_1<= rack(0);
      type_cast_2299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2299_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_1150,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv283_2300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2319_inst
    process(sext352_2316) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext352_2316(63 downto 0);
      type_cast_2319_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2324_inst
    process(ASHR_i64_i64_2323_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_2323_wire(63 downto 0);
      conv288_2325 <= tmp_var; -- 
    end process;
    type_cast_2331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2331_inst_req_0;
      type_cast_2331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2331_inst_req_1;
      type_cast_2331_inst_ack_1<= rack(0);
      type_cast_2331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_2292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv292_2332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2341_inst_req_0;
      type_cast_2341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2341_inst_req_1;
      type_cast_2341_inst_ack_1<= rack(0);
      type_cast_2341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr295_2338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv298_2342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2351_inst_req_0;
      type_cast_2351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2351_inst_req_1;
      type_cast_2351_inst_ack_1<= rack(0);
      type_cast_2351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr301_2348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_2352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2361_inst_req_0;
      type_cast_2361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2361_inst_req_1;
      type_cast_2361_inst_ack_1<= rack(0);
      type_cast_2361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr307_2358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv310_2362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2371_inst_req_0;
      type_cast_2371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2371_inst_req_1;
      type_cast_2371_inst_ack_1<= rack(0);
      type_cast_2371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr313_2368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv316_2372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2381_inst_req_0;
      type_cast_2381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2381_inst_req_1;
      type_cast_2381_inst_ack_1<= rack(0);
      type_cast_2381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2381_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr319_2378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_2382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2391_inst_req_0;
      type_cast_2391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2391_inst_req_1;
      type_cast_2391_inst_ack_1<= rack(0);
      type_cast_2391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr325_2388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv328_2392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2401_inst_req_0;
      type_cast_2401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2401_inst_req_1;
      type_cast_2401_inst_ack_1<= rack(0);
      type_cast_2401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr331_2398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv334_2402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1370_index_1_rename
    process(R_indvar425_1369_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar425_1369_resized;
      ov(13 downto 0) := iv;
      R_indvar425_1369_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1370_index_1_resize
    process(indvar425_1358) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar425_1358;
      ov := iv(13 downto 0);
      R_indvar425_1369_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1370_root_address_inst
    process(array_obj_ref_1370_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1370_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1370_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1686_index_1_rename
    process(R_ix_x0x_xlcssa_1685_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1685_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1685_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1686_index_1_resize
    process(ix_x0x_xlcssa_1552) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1552;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1685_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1686_root_address_inst
    process(array_obj_ref_1686_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1686_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1686_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1831_index_1_rename
    process(R_indvar411_1830_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar411_1830_resized;
      ov(13 downto 0) := iv;
      R_indvar411_1830_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1831_index_1_resize
    process(indvar411_1819) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar411_1819;
      ov := iv(13 downto 0);
      R_indvar411_1830_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1831_root_address_inst
    process(array_obj_ref_1831_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1831_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1831_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2151_index_1_rename
    process(R_ix_x1x_xlcssa_2150_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_2150_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_2150_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2151_index_1_resize
    process(ix_x1x_xlcssa_2013) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_2013;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_2150_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2151_root_address_inst
    process(array_obj_ref_2151_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2151_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2151_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1507_addr_0
    process(ptr_deref_1507_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1507_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1507_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1507_base_resize
    process(arrayidx_1372) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1372;
      ov := iv(13 downto 0);
      ptr_deref_1507_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1507_gather_scatter
    process(add132_1505) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_1505;
      ov(63 downto 0) := iv;
      ptr_deref_1507_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1507_root_address_inst
    process(ptr_deref_1507_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1507_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1507_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_addr_0
    process(ptr_deref_1690_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1690_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1690_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_base_resize
    process(arrayidx143_1688) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1688;
      ov := iv(13 downto 0);
      ptr_deref_1690_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_gather_scatter
    process(shl14x_xi_1681) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1681;
      ov(63 downto 0) := iv;
      ptr_deref_1690_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_root_address_inst
    process(ptr_deref_1690_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1690_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1690_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1968_addr_0
    process(ptr_deref_1968_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1968_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1968_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1968_base_resize
    process(arrayidx211_1833) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1833;
      ov := iv(13 downto 0);
      ptr_deref_1968_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1968_gather_scatter
    process(add207_1966) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_1966;
      ov(63 downto 0) := iv;
      ptr_deref_1968_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1968_root_address_inst
    process(ptr_deref_1968_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1968_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1968_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2155_addr_0
    process(ptr_deref_2155_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2155_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2155_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2155_base_resize
    process(arrayidx226_2153) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_2153;
      ov := iv(13 downto 0);
      ptr_deref_2155_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2155_gather_scatter
    process(shl14x_xi372_2146) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi372_2146;
      ov(63 downto 0) := iv;
      ptr_deref_2155_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2155_root_address_inst
    process(ptr_deref_2155_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2155_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2155_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_addr_0
    process(ptr_deref_2169_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2169_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2169_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_base_resize
    process(iNsTr_48_2167) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_48_2167;
      ov := iv(13 downto 0);
      ptr_deref_2169_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_gather_scatter
    process(type_cast_2171_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2171_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2169_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_root_address_inst
    process(ptr_deref_2169_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2169_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2169_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1280_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp383_1279;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1280_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1280_branch_req_0,
          ack0 => if_stmt_1280_branch_ack_0,
          ack1 => if_stmt_1280_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1521_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond28_1520;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1521_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1521_branch_req_0,
          ack0 => if_stmt_1521_branch_ack_0,
          ack1 => if_stmt_1521_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1572_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1571;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1572_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1572_branch_req_0,
          ack0 => if_stmt_1572_branch_ack_0,
          ack1 => if_stmt_1572_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1647_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1646;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1647_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1647_branch_req_0,
          ack0 => if_stmt_1647_branch_ack_0,
          ack1 => if_stmt_1647_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1743_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161379_1742;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1743_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1743_branch_req_0,
          ack0 => if_stmt_1743_branch_ack_0,
          ack1 => if_stmt_1743_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1982_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1981;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1982_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1982_branch_req_0,
          ack0 => if_stmt_1982_branch_ack_0,
          ack1 => if_stmt_1982_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2033_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_2032;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2033_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2033_branch_req_0,
          ack0 => if_stmt_2033_branch_ack_0,
          ack1 => if_stmt_2033_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2112_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi364_2111;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2112_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2112_branch_req_0,
          ack0 => if_stmt_2112_branch_ack_0,
          ack1 => if_stmt_2112_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2261_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_2260;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2261_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2261_branch_req_0,
          ack0 => if_stmt_2261_branch_ack_0,
          ack1 => if_stmt_2261_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1612_inst
    process(nx_x022x_xi_1593) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_1593, type_cast_1611_wire_constant, tmp_var);
      tmp_1613 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1618_inst
    process(nx_x022x_xi_1593) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_1593, type_cast_1617_wire_constant, tmp_var);
      iNsTr_35_1619 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2077_inst
    process(nx_x022x_xi357_2058) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_2058, type_cast_2076_wire_constant, tmp_var);
      tmp388_2078 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2083_inst
    process(nx_x022x_xi357_2058) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_2058, type_cast_2082_wire_constant, tmp_var);
      iNsTr_71_2084 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2190_inst
    process(add53_1200) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_1200, type_cast_2189_wire_constant, tmp_var);
      tmp389_2191 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1514_inst
    process(indvar425_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar425_1358, type_cast_1513_wire_constant, tmp_var);
      indvarx_xnext426_1515 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1975_inst
    process(indvar411_1819) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar411_1819, type_cast_1974_wire_constant, tmp_var);
      indvarx_xnext412_1976 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2205_inst
    process(tmp3_2200) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2200, type_cast_2204_wire_constant, tmp_var);
      tmp4_2206 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2254_inst
    process(indvar_2218) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2218, type_cast_2253_wire_constant, tmp_var);
      indvarx_xnext_2255 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1589_inst
    process(conv2x_xi_1584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_1584, type_cast_1588_wire_constant, tmp_var);
      shlx_xi_1590 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2054_inst
    process(conv2x_xi354_2049) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi354_2049, type_cast_2053_wire_constant, tmp_var);
      shlx_xi355_2055 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1564_inst
    process(conv83_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_1273, type_cast_1563_wire_constant, tmp_var);
      and_1565 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1669_inst
    process(Bx_xnot_1664) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1664, type_cast_1668_wire_constant, tmp_var);
      add1216x_xi_1670 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2025_inst
    process(conv155_1736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1736, type_cast_2024_wire_constant, tmp_var);
      and217_2026 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2134_inst
    process(iNsTr_97_2129) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_97_2129, type_cast_2133_wire_constant, tmp_var);
      add1216x_xi370_2135 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2241_inst
    process(mul253_2230) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul253_2230, type_cast_2240_wire_constant, tmp_var);
      conv254_2242 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1547_inst
    process(type_cast_1543_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1543_wire, type_cast_1546_wire_constant, tmp_var);
      ASHR_i64_i64_1547_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1734_inst
    process(type_cast_1730_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1730_wire, type_cast_1733_wire_constant, tmp_var);
      ASHR_i64_i64_1734_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_2008_inst
    process(type_cast_2004_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2004_wire, type_cast_2007_wire_constant, tmp_var);
      ASHR_i64_i64_2008_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_2323_inst
    process(type_cast_2319_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2319_wire, type_cast_2322_wire_constant, tmp_var);
      ASHR_i64_i64_2323_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1519_inst
    process(indvarx_xnext426_1515, umax27_1355) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext426_1515, umax27_1355, tmp_var);
      exitcond28_1520 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1570_inst
    process(and_1565) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_1565, type_cast_1569_wire_constant, tmp_var);
      tobool_1571 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1980_inst
    process(indvarx_xnext412_1976, umax19_1816) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext412_1976, umax19_1816, tmp_var);
      exitcond_1981 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2031_inst
    process(and217_2026) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_2026, type_cast_2030_wire_constant, tmp_var);
      tobool218_2032 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2259_inst
    process(indvarx_xnext_2255, tmp4_2206) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_2255, tmp4_2206, tmp_var);
      exitcond5_2260 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1306_inst
    process(tmp418_1301) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp418_1301, type_cast_1305_wire_constant, tmp_var);
      tmp419_1307 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1341_inst
    process(tmp24_1336) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp24_1336, type_cast_1340_wire_constant, tmp_var);
      tmp25_1342 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1754_inst
    process(conv155_1736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1736, type_cast_1753_wire_constant, tmp_var);
      tmp406_1755 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1802_inst
    process(tmp16_1797) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp16_1797, type_cast_1801_wire_constant, tmp_var);
      tmp17_1803 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2337_inst
    process(sub_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2292, type_cast_2336_wire_constant, tmp_var);
      shr295_2338 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2347_inst
    process(sub_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2292, type_cast_2346_wire_constant, tmp_var);
      shr301_2348 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2357_inst
    process(sub_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2292, type_cast_2356_wire_constant, tmp_var);
      shr307_2358 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2367_inst
    process(sub_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2292, type_cast_2366_wire_constant, tmp_var);
      shr313_2368 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2377_inst
    process(sub_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2292, type_cast_2376_wire_constant, tmp_var);
      shr319_2378 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2387_inst
    process(sub_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2292, type_cast_2386_wire_constant, tmp_var);
      shr325_2388 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2397_inst
    process(sub_2292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2292, type_cast_2396_wire_constant, tmp_var);
      shr331_2398 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2195_inst
    process(add73_1250, add23_1125) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1250, add23_1125, tmp_var);
      tmp393_2196 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1262_inst
    process(conv79_1254, add_1075) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_1254, add_1075, tmp_var);
      mul_1263 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1267_inst
    process(mul_1263, conv81_1258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1263, conv81_1258, tmp_var);
      mul82_1268 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1290_inst
    process(add_1075, conv79_1254) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1075, conv79_1254, tmp_var);
      tmp415_1291 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1295_inst
    process(tmp415_1291, conv81_1258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp415_1291, conv81_1258, tmp_var);
      tmp417_1296 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1321_inst
    process(add_1075, tmp20_1317) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1075, tmp20_1317, tmp_var);
      tmp21_1322 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1330_inst
    process(tmp21_1322, tmp22_1326) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp21_1322, tmp22_1326, tmp_var);
      tmp23_1331 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1710_inst
    process(conv153_1706, conv145_1698) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1706, conv145_1698, tmp_var);
      mul148_1711 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1715_inst
    process(mul148_1711, add63_1225) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1711, add63_1225, tmp_var);
      mul151_1716 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1720_inst
    process(mul151_1716, conv147_1702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1716, conv147_1702, tmp_var);
      mul154_1721 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1769_inst
    process(add63_1225, tmp9_1765) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_1225, tmp9_1765, tmp_var);
      tmp10_1770 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1778_inst
    process(tmp10_1770, tmp11_1774) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp10_1770, tmp11_1774, tmp_var);
      tmp12_1779 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1787_inst
    process(tmp12_1779, tmp13_1783) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1779, tmp13_1783, tmp_var);
      tmp14_1788 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2214_inst
    process(add63_1225, tmp6_2210) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_1225, tmp6_2210, tmp_var);
      tmp7_2215 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2229_inst
    process(tmp7_2215, indvar_2218) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp7_2215, indvar_2218, tmp_var);
      mul253_2230 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2310_inst
    process(mul284_2306, conv281_2296) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul284_2306, conv281_2296, tmp_var);
      mul287_2311 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2315_inst
    process(mul287_2311, conv153_1706) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul287_2311, conv153_1706, tmp_var);
      sext352_2316 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1099_inst
    process(shl10_1088, conv12_1095) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_1088, conv12_1095, tmp_var);
      add13_1100 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1124_inst
    process(shl20_1113, conv22_1120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_1113, conv22_1120, tmp_var);
      add23_1125 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1149_inst
    process(shl30_1138, conv32_1145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_1138, conv32_1145, tmp_var);
      add33_1150 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1174_inst
    process(shl40_1163, conv42_1170) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_1163, conv42_1170, tmp_var);
      add43_1175 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1199_inst
    process(shl50_1188, conv52_1195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_1188, conv52_1195, tmp_var);
      add53_1200 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1249_inst
    process(shl70_1238, conv72_1245) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_1238, conv72_1245, tmp_var);
      add73_1250 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1074_inst
    process(shl_1063, conv3_1070) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1063, conv3_1070, tmp_var);
      add_1075 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1224_inst
    process(shl60_1213, conv62_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_1213, conv62_1220, tmp_var);
      add63_1225 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1396_inst
    process(shl92_1385, conv95_1392) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_1385, conv95_1392, tmp_var);
      add96_1397 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1414_inst
    process(shl98_1403, conv101_1410) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_1403, conv101_1410, tmp_var);
      add102_1415 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1432_inst
    process(shl104_1421, conv107_1428) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_1421, conv107_1428, tmp_var);
      add108_1433 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1450_inst
    process(shl110_1439, conv113_1446) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_1439, conv113_1446, tmp_var);
      add114_1451 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1468_inst
    process(shl116_1457, conv119_1464) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_1457, conv119_1464, tmp_var);
      add120_1469 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1486_inst
    process(shl122_1475, conv125_1482) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_1475, conv125_1482, tmp_var);
      add126_1487 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1504_inst
    process(shl128_1493, conv131_1500) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_1493, conv131_1500, tmp_var);
      add132_1505 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1630_inst
    process(conv5x_xi_1626, elementx_x021x_xi_1600) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1626, elementx_x021x_xi_1600, tmp_var);
      addx_xi_1631 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1857_inst
    process(shl167_1846, conv170_1853) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1846, conv170_1853, tmp_var);
      add171_1858 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1875_inst
    process(shl173_1864, conv176_1871) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1864, conv176_1871, tmp_var);
      add177_1876 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1893_inst
    process(shl179_1882, conv182_1889) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1882, conv182_1889, tmp_var);
      add183_1894 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1911_inst
    process(shl185_1900, conv188_1907) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1900, conv188_1907, tmp_var);
      add189_1912 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1929_inst
    process(shl191_1918, conv194_1925) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1918, conv194_1925, tmp_var);
      add195_1930 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1947_inst
    process(shl197_1936, conv200_1943) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_1936, conv200_1943, tmp_var);
      add201_1948 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1965_inst
    process(shl203_1954, conv206_1961) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_1954, conv206_1961, tmp_var);
      add207_1966 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2095_inst
    process(conv5x_xi360_2091, elementx_x021x_xi358_2065) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi360_2091, elementx_x021x_xi358_2065, tmp_var);
      addx_xi361_2096 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1087_inst
    process(conv9_1082) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_1082, type_cast_1086_wire_constant, tmp_var);
      shl10_1088 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1112_inst
    process(conv19_1107) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_1107, type_cast_1111_wire_constant, tmp_var);
      shl20_1113 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1137_inst
    process(conv29_1132) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_1132, type_cast_1136_wire_constant, tmp_var);
      shl30_1138 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1162_inst
    process(conv39_1157) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_1157, type_cast_1161_wire_constant, tmp_var);
      shl40_1163 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1187_inst
    process(conv49_1182) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1182, type_cast_1186_wire_constant, tmp_var);
      shl50_1188 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1237_inst
    process(conv69_1232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_1232, type_cast_1236_wire_constant, tmp_var);
      shl70_1238 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1062_inst
    process(conv1_1057) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_1057, type_cast_1061_wire_constant, tmp_var);
      shl_1063 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1583_inst
    process(mul82_1268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_1268, type_cast_1582_wire_constant, tmp_var);
      conv2x_xi_1584 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1212_inst
    process(conv59_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_1207, type_cast_1211_wire_constant, tmp_var);
      shl60_1213 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1384_inst
    process(conv90_1379) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_1379, type_cast_1383_wire_constant, tmp_var);
      shl92_1385 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1402_inst
    process(add96_1397) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_1397, type_cast_1401_wire_constant, tmp_var);
      shl98_1403 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1420_inst
    process(add102_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_1415, type_cast_1419_wire_constant, tmp_var);
      shl104_1421 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1438_inst
    process(add108_1433) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_1433, type_cast_1437_wire_constant, tmp_var);
      shl110_1439 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1456_inst
    process(add114_1451) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_1451, type_cast_1455_wire_constant, tmp_var);
      shl116_1457 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1474_inst
    process(add120_1469) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_1469, type_cast_1473_wire_constant, tmp_var);
      shl122_1475 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1492_inst
    process(add126_1487) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_1487, type_cast_1491_wire_constant, tmp_var);
      shl128_1493 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1539_inst
    process(umax421_1534) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax421_1534, type_cast_1538_wire_constant, tmp_var);
      tmp422_1540 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1636_inst
    process(addx_xi_1631) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1631, type_cast_1635_wire_constant, tmp_var);
      shl8x_xi_1637 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1663_inst
    process(conv83_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_1273, type_cast_1662_wire_constant, tmp_var);
      Bx_xnot_1664 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1680_inst
    process(shl8x_xix_xlcssa_1654, sh_promx_xi_1676) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1654, sh_promx_xi_1676, tmp_var);
      shl14x_xi_1681 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1726_inst
    process(mul154_1721) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1721, type_cast_1725_wire_constant, tmp_var);
      sext_1727 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1845_inst
    process(conv165_1840) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1840, type_cast_1844_wire_constant, tmp_var);
      shl167_1846 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1863_inst
    process(add171_1858) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1858, type_cast_1862_wire_constant, tmp_var);
      shl173_1864 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1881_inst
    process(add177_1876) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1876, type_cast_1880_wire_constant, tmp_var);
      shl179_1882 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1899_inst
    process(add183_1894) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1894, type_cast_1898_wire_constant, tmp_var);
      shl185_1900 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1917_inst
    process(add189_1912) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1912, type_cast_1916_wire_constant, tmp_var);
      shl191_1918 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1935_inst
    process(add195_1930) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_1930, type_cast_1934_wire_constant, tmp_var);
      shl197_1936 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1953_inst
    process(add201_1948) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_1948, type_cast_1952_wire_constant, tmp_var);
      shl203_1954 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2000_inst
    process(umax_1995) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1995, type_cast_1999_wire_constant, tmp_var);
      tmp408_2001 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2044_inst
    process(mul154_1721) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1721, type_cast_2043_wire_constant, tmp_var);
      iNsTr_59_2045 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2101_inst
    process(addx_xi361_2096) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi361_2096, type_cast_2100_wire_constant, tmp_var);
      shl8x_xi362_2102 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2128_inst
    process(mul154_1721) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1721, type_cast_2127_wire_constant, tmp_var);
      iNsTr_97_2129 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2145_inst
    process(shl8x_xi362x_xlcssa_2119, sh_promx_xi371_2141) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi362x_xlcssa_2119, sh_promx_xi371_2141, tmp_var);
      shl14x_xi372_2146 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2305_inst
    process(conv283_2300) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv283_2300, type_cast_2304_wire_constant, tmp_var);
      mul284_2306 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_2291_inst
    process(conv276_2287, conv230_2272) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv276_2287, conv230_2272, tmp_var);
      sub_2292 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1278_inst
    process(mul82_1268) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_1268, type_cast_1277_wire_constant, tmp_var);
      cmp383_1279 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1312_inst
    process(tmp419_1307) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp419_1307, type_cast_1311_wire_constant, tmp_var);
      tmp420_1313 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1347_inst
    process(tmp25_1342) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp25_1342, type_cast_1346_wire_constant, tmp_var);
      tmp26_1348 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1741_inst
    process(conv155_1736) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1736, type_cast_1740_wire_constant, tmp_var);
      cmp161379_1742 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1760_inst
    process(tmp406_1755) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp406_1755, type_cast_1759_wire_constant, tmp_var);
      tmp407_1761 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1808_inst
    process(tmp17_1803) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp17_1803, type_cast_1807_wire_constant, tmp_var);
      tmp18_1809 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1645_inst
    process(convx_xi_1641, shlx_xi_1590) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1641, shlx_xi_1590, tmp_var);
      cmpx_xi_1646 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2110_inst
    process(convx_xi363_2106, shlx_xi355_2055) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi363_2106, shlx_xi355_2055, tmp_var);
      cmpx_xi364_2111 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1675_inst
    process(add1216x_xi_1670) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1670, type_cast_1674_wire_constant, tmp_var);
      sh_promx_xi_1676 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_2140_inst
    process(add1216x_xi370_2135) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi370_2135, type_cast_2139_wire_constant, tmp_var);
      sh_promx_xi371_2141 <= tmp_var; --
    end process;
    -- shared split operator group (122) : array_obj_ref_1370_index_offset 
    ApIntAdd_group_122: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar425_1369_scaled;
      array_obj_ref_1370_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1370_index_offset_req_0;
      array_obj_ref_1370_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1370_index_offset_req_1;
      array_obj_ref_1370_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_122_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_122_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : array_obj_ref_1686_index_offset 
    ApIntAdd_group_123: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1685_scaled;
      array_obj_ref_1686_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1686_index_offset_req_0;
      array_obj_ref_1686_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1686_index_offset_req_1;
      array_obj_ref_1686_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_123_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_123_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : array_obj_ref_1831_index_offset 
    ApIntAdd_group_124: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar411_1830_scaled;
      array_obj_ref_1831_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1831_index_offset_req_0;
      array_obj_ref_1831_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1831_index_offset_req_1;
      array_obj_ref_1831_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_124_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_124_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : array_obj_ref_2151_index_offset 
    ApIntAdd_group_125: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_2150_scaled;
      array_obj_ref_2151_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2151_index_offset_req_0;
      array_obj_ref_2151_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2151_index_offset_req_1;
      array_obj_ref_2151_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_125_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_125_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- unary operator type_cast_1271_inst
    process(mul82_1268) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_1268, tmp_var);
      type_cast_1271_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1299_inst
    process(tmp417_1296) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp417_1296, tmp_var);
      type_cast_1299_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1334_inst
    process(tmp23_1331) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp23_1331, tmp_var);
      type_cast_1334_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1795_inst
    process(tmp15_1792) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp15_1792, tmp_var);
      type_cast_1795_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2270_inst
    process(call229_2175) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_2175, tmp_var);
      type_cast_2270_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2285_inst
    process(call275_2282) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_2282, tmp_var);
      type_cast_2285_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1690_store_0 ptr_deref_1507_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1690_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1507_store_0_req_0;
      ptr_deref_1690_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1507_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1690_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1507_store_0_req_1;
      ptr_deref_1690_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1507_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1690_word_address_0 & ptr_deref_1507_word_address_0;
      data_in <= ptr_deref_1690_data_0 & ptr_deref_1507_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1968_store_0 ptr_deref_2155_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1968_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2155_store_0_req_0;
      ptr_deref_1968_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2155_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1968_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2155_store_0_req_1;
      ptr_deref_1968_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2155_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1968_word_address_0 & ptr_deref_2155_word_address_0;
      data_in <= ptr_deref_1968_data_0 & ptr_deref_2155_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_2169_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2169_store_0_req_0;
      ptr_deref_2169_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2169_store_0_req_1;
      ptr_deref_2169_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2169_word_address_0;
      data_in <= ptr_deref_2169_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_input_done_pipe_2274_inst RPIPE_input_done_pipe_2278_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_input_done_pipe_2274_inst_req_0;
      reqL_unguarded(0) <= RPIPE_input_done_pipe_2278_inst_req_0;
      RPIPE_input_done_pipe_2274_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_input_done_pipe_2278_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_input_done_pipe_2274_inst_req_1;
      reqR_unguarded(0) <= RPIPE_input_done_pipe_2278_inst_req_1;
      RPIPE_input_done_pipe_2274_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_input_done_pipe_2278_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      call270_2275 <= data_out(15 downto 8);
      call273_2279 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_maxpool_input_pipe_1848_inst RPIPE_maxpool_input_pipe_1866_inst RPIPE_maxpool_input_pipe_1884_inst RPIPE_maxpool_input_pipe_1902_inst RPIPE_maxpool_input_pipe_1920_inst RPIPE_maxpool_input_pipe_1938_inst RPIPE_maxpool_input_pipe_1835_inst RPIPE_maxpool_input_pipe_1052_inst RPIPE_maxpool_input_pipe_1065_inst RPIPE_maxpool_input_pipe_1077_inst RPIPE_maxpool_input_pipe_1090_inst RPIPE_maxpool_input_pipe_1102_inst RPIPE_maxpool_input_pipe_1115_inst RPIPE_maxpool_input_pipe_1127_inst RPIPE_maxpool_input_pipe_1140_inst RPIPE_maxpool_input_pipe_1152_inst RPIPE_maxpool_input_pipe_1165_inst RPIPE_maxpool_input_pipe_1177_inst RPIPE_maxpool_input_pipe_1190_inst RPIPE_maxpool_input_pipe_1202_inst RPIPE_maxpool_input_pipe_1215_inst RPIPE_maxpool_input_pipe_1227_inst RPIPE_maxpool_input_pipe_1240_inst RPIPE_maxpool_input_pipe_1374_inst RPIPE_maxpool_input_pipe_1387_inst RPIPE_maxpool_input_pipe_1405_inst RPIPE_maxpool_input_pipe_1423_inst RPIPE_maxpool_input_pipe_1441_inst RPIPE_maxpool_input_pipe_1459_inst RPIPE_maxpool_input_pipe_1477_inst RPIPE_maxpool_input_pipe_1495_inst RPIPE_maxpool_input_pipe_1621_inst RPIPE_maxpool_input_pipe_1956_inst RPIPE_maxpool_input_pipe_2086_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_1848_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_1866_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_1884_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_1902_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_1920_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_1938_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_1835_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_1052_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_1065_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_1077_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_1090_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_1102_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_1115_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_1127_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1140_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_1152_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_1165_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_1177_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_1190_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_1202_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_1215_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_1227_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1240_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1374_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1387_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1405_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1423_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1441_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1459_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1477_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1495_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1621_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1956_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_2086_inst_req_0;
      RPIPE_maxpool_input_pipe_1848_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_1866_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_1884_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_1902_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_1920_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_1938_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_1835_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_1052_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_1065_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_1077_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_1090_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_1102_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_1115_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_1127_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1140_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_1152_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_1165_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_1177_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_1190_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_1202_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_1215_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_1227_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_1240_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1374_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1387_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1405_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1423_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1441_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1459_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1477_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1495_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1621_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1956_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_2086_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_1848_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_1866_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_1884_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_1902_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_1920_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_1938_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_1835_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_1052_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_1065_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_1077_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_1090_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_1102_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_1115_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_1127_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1140_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_1152_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_1165_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_1177_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_1190_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_1202_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_1215_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_1227_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1240_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1374_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1387_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1405_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1423_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1441_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1459_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1477_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1495_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1621_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1956_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_2086_inst_req_1;
      RPIPE_maxpool_input_pipe_1848_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_1866_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_1884_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_1902_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_1920_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_1938_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_1835_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_1052_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_1065_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_1077_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_1090_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_1102_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_1115_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_1127_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1140_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_1152_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_1165_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_1177_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_1190_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_1202_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_1215_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_1227_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_1240_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1374_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1387_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1405_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1423_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1441_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1459_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1477_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1495_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1621_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1956_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_2086_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call168_1849 <= data_out(271 downto 264);
      call174_1867 <= data_out(263 downto 256);
      call180_1885 <= data_out(255 downto 248);
      call186_1903 <= data_out(247 downto 240);
      call192_1921 <= data_out(239 downto 232);
      call198_1939 <= data_out(231 downto 224);
      call164_1836 <= data_out(223 downto 216);
      call_1053 <= data_out(215 downto 208);
      call2_1066 <= data_out(207 downto 200);
      call6_1078 <= data_out(199 downto 192);
      call11_1091 <= data_out(191 downto 184);
      call16_1103 <= data_out(183 downto 176);
      call21_1116 <= data_out(175 downto 168);
      call26_1128 <= data_out(167 downto 160);
      call31_1141 <= data_out(159 downto 152);
      call36_1153 <= data_out(151 downto 144);
      call41_1166 <= data_out(143 downto 136);
      call46_1178 <= data_out(135 downto 128);
      call51_1191 <= data_out(127 downto 120);
      call56_1203 <= data_out(119 downto 112);
      call61_1216 <= data_out(111 downto 104);
      call66_1228 <= data_out(103 downto 96);
      call71_1241 <= data_out(95 downto 88);
      call89_1375 <= data_out(87 downto 80);
      call93_1388 <= data_out(79 downto 72);
      call99_1406 <= data_out(71 downto 64);
      call105_1424 <= data_out(63 downto 56);
      call111_1442 <= data_out(55 downto 48);
      call117_1460 <= data_out(47 downto 40);
      call123_1478 <= data_out(39 downto 32);
      call129_1496 <= data_out(31 downto 24);
      callx_xi_1622 <= data_out(23 downto 16);
      call204_1957 <= data_out(15 downto 8);
      callx_xi359_2087 <= data_out(7 downto 0);
      maxpool_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_1_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_1", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_2403_inst WPIPE_maxpool_output_pipe_2406_inst WPIPE_maxpool_output_pipe_2409_inst WPIPE_maxpool_output_pipe_2412_inst WPIPE_maxpool_output_pipe_2415_inst WPIPE_maxpool_output_pipe_2418_inst WPIPE_maxpool_output_pipe_2421_inst WPIPE_maxpool_output_pipe_2424_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2403_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2406_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2409_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2412_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2415_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2418_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2421_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2424_inst_req_0;
      WPIPE_maxpool_output_pipe_2403_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2406_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2409_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2412_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2415_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2418_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2421_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2424_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2403_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2406_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2409_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2412_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2415_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2418_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2421_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2424_inst_req_1;
      WPIPE_maxpool_output_pipe_2403_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2406_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2409_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2412_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2415_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2418_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2421_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2424_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv334_2402 & conv328_2392 & conv322_2382 & conv316_2372 & conv310_2362 & conv304_2352 & conv298_2342 & conv292_2332;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_2231_inst WPIPE_num_out_pipe_2234_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_num_out_pipe_2231_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_2234_inst_req_0;
      WPIPE_num_out_pipe_2231_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_num_out_pipe_2234_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_num_out_pipe_2231_inst_req_1;
      update_req_unguarded(0) <= WPIPE_num_out_pipe_2234_inst_req_1;
      WPIPE_num_out_pipe_2231_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_num_out_pipe_2234_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= add33_1150 & add43_1175;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_output_pipe_2176_inst WPIPE_output_pipe_2179_inst WPIPE_output_pipe_2182_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal sample_req, sample_ack : BooleanArray( 2 downto 0);
      signal update_req, update_ack : BooleanArray( 2 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 2 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      sample_req_unguarded(2) <= WPIPE_output_pipe_2176_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_output_pipe_2179_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_output_pipe_2182_inst_req_0;
      WPIPE_output_pipe_2176_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_output_pipe_2179_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_output_pipe_2182_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(2) <= WPIPE_output_pipe_2176_inst_req_1;
      update_req_unguarded(1) <= WPIPE_output_pipe_2179_inst_req_1;
      update_req_unguarded(0) <= WPIPE_output_pipe_2182_inst_req_1;
      WPIPE_output_pipe_2176_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_output_pipe_2179_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_output_pipe_2182_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      data_in <= add33_1150 & add43_1175 & add53_1200;
      output_pipe_write_2_gI: SplitGuardInterface generic map(name => "output_pipe_write_2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 3, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_2175_call call_stmt_2282_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2175_call_req_0;
      reqL_unguarded(0) <= call_stmt_2282_call_req_0;
      call_stmt_2175_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2282_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2175_call_req_1;
      reqR_unguarded(0) <= call_stmt_2282_call_req_1;
      call_stmt_2175_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2282_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_2175 <= data_out(127 downto 64);
      call275_2282 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2245_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2245_call_req_0;
      call_stmt_2245_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2245_call_req_1;
      call_stmt_2245_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv254_2242 & add23_1125;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(79 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2249_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2249_call_req_0;
      call_stmt_2249_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2249_call_req_1;
      call_stmt_2249_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add33_1150 & add23_1125 & add13_1100;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(47 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_2327_call 
    sendB_call_group_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2327_call_req_0;
      call_stmt_2327_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2327_call_req_1;
      call_stmt_2327_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv288_2325;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(63 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_6200_start: Boolean;
  signal convolve_CP_6200_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_xxconvolvexxconv_k2_2738_inst_ack_1 : boolean;
  signal type_cast_2801_inst_ack_0 : boolean;
  signal do_while_stmt_2455_branch_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2738_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2745_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2745_inst_req_1 : boolean;
  signal W_num_done_2703_delayed_1_0_2786_inst_req_0 : boolean;
  signal W_store_kernel_2660_delayed_1_0_2741_inst_ack_0 : boolean;
  signal W_num_done_2703_delayed_1_0_2786_inst_ack_0 : boolean;
  signal type_cast_2801_inst_req_1 : boolean;
  signal W_store_kernel_2660_delayed_1_0_2741_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2799_inst_req_0 : boolean;
  signal W_store_kernel_2660_delayed_1_0_2741_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_2806_inst_ack_1 : boolean;
  signal n_col_2777_2472_buf_req_1 : boolean;
  signal n_col_2777_2472_buf_ack_1 : boolean;
  signal n_row_2785_2467_buf_req_0 : boolean;
  signal n_chl_2755_2483_buf_req_0 : boolean;
  signal n_chl_2755_2483_buf_ack_0 : boolean;
  signal n_row_2785_2467_buf_ack_1 : boolean;
  signal phi_stmt_2479_ack_0 : boolean;
  signal n_row_2785_2467_buf_ack_0 : boolean;
  signal W_num_done_2708_delayed_1_0_2795_inst_req_1 : boolean;
  signal phi_stmt_2468_ack_0 : boolean;
  signal n_num_2766_2478_buf_req_1 : boolean;
  signal W_num_done_2708_delayed_1_0_2795_inst_ack_1 : boolean;
  signal phi_stmt_2468_req_1 : boolean;
  signal phi_stmt_2473_req_1 : boolean;
  signal n_col_2777_2472_buf_ack_0 : boolean;
  signal phi_stmt_2468_req_0 : boolean;
  signal n_num_2766_2478_buf_ack_1 : boolean;
  signal phi_stmt_2473_req_0 : boolean;
  signal phi_stmt_2473_ack_0 : boolean;
  signal n_num_2766_2478_buf_req_0 : boolean;
  signal n_chl_2755_2483_buf_req_1 : boolean;
  signal W_num_done_2708_delayed_1_0_2795_inst_ack_0 : boolean;
  signal n_chl_2755_2483_buf_ack_1 : boolean;
  signal WPIPE_output_pipe_2799_inst_ack_0 : boolean;
  signal phi_stmt_2479_req_0 : boolean;
  signal n_num_2766_2478_buf_ack_0 : boolean;
  signal n_row_2785_2467_buf_req_1 : boolean;
  signal phi_stmt_2479_req_1 : boolean;
  signal do_while_stmt_2455_branch_ack_1 : boolean;
  signal W_store_kernel_2660_delayed_1_0_2741_inst_ack_1 : boolean;
  signal W_num_done_2703_delayed_1_0_2786_inst_req_1 : boolean;
  signal type_cast_2801_inst_req_0 : boolean;
  signal type_cast_2801_inst_ack_1 : boolean;
  signal W_num_done_2703_delayed_1_0_2786_inst_ack_1 : boolean;
  signal W_store_kernel_2656_delayed_1_0_2734_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2738_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_2806_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2441_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2441_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2441_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_2441_inst_ack_1 : boolean;
  signal SUB_u16_u16_2443_inst_req_0 : boolean;
  signal SUB_u16_u16_2443_inst_ack_0 : boolean;
  signal SUB_u16_u16_2443_inst_req_1 : boolean;
  signal SUB_u16_u16_2443_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_2446_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2446_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2446_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_2446_inst_ack_1 : boolean;
  signal SUB_u16_u16_2448_inst_req_0 : boolean;
  signal SUB_u16_u16_2448_inst_ack_0 : boolean;
  signal SUB_u16_u16_2448_inst_req_1 : boolean;
  signal SUB_u16_u16_2448_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_2451_inst_req_0 : boolean;
  signal RPIPE_size_pipe_2451_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_2451_inst_req_1 : boolean;
  signal RPIPE_size_pipe_2451_inst_ack_1 : boolean;
  signal SUB_u16_u16_2453_inst_req_0 : boolean;
  signal SUB_u16_u16_2453_inst_ack_0 : boolean;
  signal SUB_u16_u16_2453_inst_req_1 : boolean;
  signal SUB_u16_u16_2453_inst_ack_1 : boolean;
  signal do_while_stmt_2455_branch_req_0 : boolean;
  signal phi_stmt_2457_req_1 : boolean;
  signal phi_stmt_2457_req_0 : boolean;
  signal phi_stmt_2457_ack_0 : boolean;
  signal n_col_2777_2472_buf_req_0 : boolean;
  signal nacc_2794_2462_buf_req_0 : boolean;
  signal nacc_2794_2462_buf_ack_0 : boolean;
  signal nacc_2794_2462_buf_req_1 : boolean;
  signal nacc_2794_2462_buf_ack_1 : boolean;
  signal phi_stmt_2463_req_1 : boolean;
  signal phi_stmt_2463_req_0 : boolean;
  signal phi_stmt_2463_ack_0 : boolean;
  signal RPIPE_input_pipe1_2496_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_2496_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_2496_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_2496_inst_ack_1 : boolean;
  signal RPIPE_input_pipe2_2500_inst_req_0 : boolean;
  signal RPIPE_input_pipe2_2500_inst_ack_0 : boolean;
  signal RPIPE_input_pipe2_2500_inst_req_1 : boolean;
  signal RPIPE_input_pipe2_2500_inst_ack_1 : boolean;
  signal W_store_kernel_2656_delayed_1_0_2734_inst_ack_1 : boolean;
  signal W_store_kernel_2656_delayed_1_0_2734_inst_req_1 : boolean;
  signal W_num_done_2708_delayed_1_0_2795_inst_req_0 : boolean;
  signal W_store_kernel_2656_delayed_1_0_2734_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_2806_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_2504_inst_req_0 : boolean;
  signal RPIPE_input_pipe3_2504_inst_ack_0 : boolean;
  signal RPIPE_input_pipe3_2504_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_2504_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2745_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2745_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2508_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2508_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2738_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2508_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2508_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2799_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2799_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_2806_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2512_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2512_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2512_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2512_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2516_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2516_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2516_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2516_inst_ack_1 : boolean;
  signal W_read_ip_2474_delayed_1_0_2518_inst_req_0 : boolean;
  signal W_read_ip_2474_delayed_1_0_2518_inst_ack_0 : boolean;
  signal W_read_ip_2474_delayed_1_0_2518_inst_req_1 : boolean;
  signal W_read_ip_2474_delayed_1_0_2518_inst_ack_1 : boolean;
  signal W_read_ip_2480_delayed_1_0_2527_inst_req_0 : boolean;
  signal W_read_ip_2480_delayed_1_0_2527_inst_ack_0 : boolean;
  signal W_read_ip_2480_delayed_1_0_2527_inst_req_1 : boolean;
  signal W_read_ip_2480_delayed_1_0_2527_inst_ack_1 : boolean;
  signal W_read_ip_2486_delayed_1_0_2536_inst_req_0 : boolean;
  signal W_read_ip_2486_delayed_1_0_2536_inst_ack_0 : boolean;
  signal W_read_ip_2486_delayed_1_0_2536_inst_req_1 : boolean;
  signal W_read_ip_2486_delayed_1_0_2536_inst_ack_1 : boolean;
  signal W_write_input_2500_delayed_1_0_2554_inst_req_0 : boolean;
  signal W_write_input_2500_delayed_1_0_2554_inst_ack_0 : boolean;
  signal W_write_input_2500_delayed_1_0_2554_inst_req_1 : boolean;
  signal W_write_input_2500_delayed_1_0_2554_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2558_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2558_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2558_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2558_inst_ack_1 : boolean;
  signal W_write_input_2504_delayed_1_0_2561_inst_req_0 : boolean;
  signal W_write_input_2504_delayed_1_0_2561_inst_ack_0 : boolean;
  signal W_write_input_2504_delayed_1_0_2561_inst_req_1 : boolean;
  signal W_write_input_2504_delayed_1_0_2561_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2565_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2565_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2565_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2565_inst_ack_1 : boolean;
  signal W_write_input_2508_delayed_1_0_2568_inst_req_0 : boolean;
  signal W_write_input_2508_delayed_1_0_2568_inst_ack_0 : boolean;
  signal W_write_input_2508_delayed_1_0_2568_inst_req_1 : boolean;
  signal W_write_input_2508_delayed_1_0_2568_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2572_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2572_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2572_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2572_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_2598_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_2598_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_2598_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_2598_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe2_2602_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_2602_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_2602_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe2_2602_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe3_2606_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe3_2606_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe3_2606_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_2606_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2610_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2610_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2610_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2610_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2614_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2614_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2614_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2614_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2618_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2618_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2618_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2618_inst_ack_1 : boolean;
  signal W_read_k_2558_delayed_1_0_2620_inst_req_0 : boolean;
  signal W_read_k_2558_delayed_1_0_2620_inst_ack_0 : boolean;
  signal W_read_k_2558_delayed_1_0_2620_inst_req_1 : boolean;
  signal W_read_k_2558_delayed_1_0_2620_inst_ack_1 : boolean;
  signal W_read_k_2564_delayed_1_0_2629_inst_req_0 : boolean;
  signal W_read_k_2564_delayed_1_0_2629_inst_ack_0 : boolean;
  signal W_read_k_2564_delayed_1_0_2629_inst_req_1 : boolean;
  signal W_read_k_2564_delayed_1_0_2629_inst_ack_1 : boolean;
  signal W_read_k_2570_delayed_1_0_2638_inst_req_0 : boolean;
  signal W_read_k_2570_delayed_1_0_2638_inst_ack_0 : boolean;
  signal W_read_k_2570_delayed_1_0_2638_inst_req_1 : boolean;
  signal W_read_k_2570_delayed_1_0_2638_inst_ack_1 : boolean;
  signal W_acc_2606_delayed_1_0_2677_inst_req_0 : boolean;
  signal W_acc_2606_delayed_1_0_2677_inst_ack_0 : boolean;
  signal W_acc_2606_delayed_1_0_2677_inst_req_1 : boolean;
  signal W_acc_2606_delayed_1_0_2677_inst_ack_1 : boolean;
  signal W_store_kernel_2652_delayed_1_0_2727_inst_req_0 : boolean;
  signal W_store_kernel_2652_delayed_1_0_2727_inst_ack_0 : boolean;
  signal W_store_kernel_2652_delayed_1_0_2727_inst_req_1 : boolean;
  signal W_store_kernel_2652_delayed_1_0_2727_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2731_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2731_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2731_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2731_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_6200_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6200_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_6200_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6200_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_6200: Block -- control-path 
    signal convolve_CP_6200_elements: BooleanArray(262 downto 0);
    -- 
  begin -- 
    convolve_CP_6200_elements(0) <= convolve_CP_6200_start;
    convolve_CP_6200_symbol <= convolve_CP_6200_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	262 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_2438/merge_stmt_2439__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_2438/merge_stmt_2439__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_2438/merge_stmt_2439_dead_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2438/$entry
      -- CP-element group 0: 	 branch_block_stmt_2438/branch_block_stmt_2438__entry__
      -- CP-element group 0: 	 branch_block_stmt_2438/merge_stmt_2439__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2438/$exit
      -- CP-element group 1: 	 branch_block_stmt_2438/branch_block_stmt_2438__exit__
      -- 
    convolve_CP_6200_elements(1) <= false; 
    -- CP-element group 2:  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	259 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	260 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2438/assign_stmt_2808/$entry
      -- CP-element group 2: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_2438/do_while_stmt_2455__exit__
      -- CP-element group 2: 	 branch_block_stmt_2438/assign_stmt_2808__entry__
      -- 
    req_7054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(2), ack => WPIPE_input_done_pipe_2806_inst_req_0); -- 
    convolve_CP_6200_elements(2) <= convolve_CP_6200_elements(259);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	262 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Update/cr
      -- 
    ra_6232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2441_inst_ack_0, ack => convolve_CP_6200_elements(3)); -- 
    cr_6236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(3), ack => RPIPE_num_out_pipe_2441_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Sample/rr
      -- 
    ca_6237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2441_inst_ack_1, ack => convolve_CP_6200_elements(4)); -- 
    rr_6241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(4), ack => SUB_u16_u16_2443_inst_req_0); -- 
    rr_6259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(4), ack => RPIPE_num_out_pipe_2446_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Sample/ra
      -- 
    ra_6242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2443_inst_ack_0, ack => convolve_CP_6200_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	262 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	15 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Update/ca
      -- 
    ca_6247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2443_inst_ack_1, ack => convolve_CP_6200_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_update_start_
      -- CP-element group 7: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Update/cr
      -- 
    ra_6260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2446_inst_ack_0, ack => convolve_CP_6200_elements(7)); -- 
    cr_6264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(7), ack => RPIPE_num_out_pipe_2446_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2446_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Sample/rr
      -- 
    ca_6265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2446_inst_ack_1, ack => convolve_CP_6200_elements(8)); -- 
    rr_6269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(8), ack => SUB_u16_u16_2448_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Sample/ra
      -- 
    ra_6270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2448_inst_ack_0, ack => convolve_CP_6200_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	262 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Update/ca
      -- 
    ca_6275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2448_inst_ack_1, ack => convolve_CP_6200_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	262 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Update/cr
      -- 
    ra_6288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2451_inst_ack_0, ack => convolve_CP_6200_elements(11)); -- 
    cr_6292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(11), ack => RPIPE_size_pipe_2451_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Sample/rr
      -- 
    ca_6293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2451_inst_ack_1, ack => convolve_CP_6200_elements(12)); -- 
    rr_6297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(12), ack => SUB_u16_u16_2453_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Sample/ra
      -- 
    ra_6298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2453_inst_ack_0, ack => convolve_CP_6200_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	262 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Update/ca
      -- 
    ca_6303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2453_inst_ack_1, ack => convolve_CP_6200_elements(14)); -- 
    -- CP-element group 15:  join  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	6 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454__exit__
      -- CP-element group 15: 	 branch_block_stmt_2438/do_while_stmt_2455__entry__
      -- CP-element group 15: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/$exit
      -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(10) & convolve_CP_6200_elements(14) & convolve_CP_6200_elements(6);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2438/do_while_stmt_2455/$entry
      -- CP-element group 16: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455__entry__
      -- 
    convolve_CP_6200_elements(16) <= convolve_CP_6200_elements(15);
    -- CP-element group 17:  merge  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	259 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455__exit__
      -- 
    -- Element group convolve_CP_6200_elements(17) is bound as output of CP function.
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_back
      -- 
    -- Element group convolve_CP_6200_elements(18) is bound as output of CP function.
    -- CP-element group 19:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	257 
    -- CP-element group 19: 	258 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_taken/$entry
      -- CP-element group 19: 	 branch_block_stmt_2438/do_while_stmt_2455/condition_done
      -- CP-element group 19: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_exit/$entry
      -- 
    convolve_CP_6200_elements(19) <= convolve_CP_6200_elements(24);
    -- CP-element group 20:  branch  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	256 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_body_done
      -- 
    convolve_CP_6200_elements(20) <= convolve_CP_6200_elements(256);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	33 
    -- CP-element group 21: 	52 
    -- CP-element group 21: 	71 
    -- CP-element group 21: 	90 
    -- CP-element group 21: 	109 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_6200_elements(21) <= convolve_CP_6200_elements(18);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	35 
    -- CP-element group 22: 	54 
    -- CP-element group 22: 	73 
    -- CP-element group 22: 	92 
    -- CP-element group 22: 	111 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_6200_elements(22) <= convolve_CP_6200_elements(16);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	255 
    -- CP-element group 23: 	29 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	47 
    -- CP-element group 23: 	66 
    -- CP-element group 23: 	84 
    -- CP-element group 23: 	65 
    -- CP-element group 23: 	85 
    -- CP-element group 23: 	103 
    -- CP-element group 23: 	104 
    -- CP-element group 23: 	126 
    -- CP-element group 23: 	122 
    -- CP-element group 23: 	130 
    -- CP-element group 23: 	134 
    -- CP-element group 23: 	138 
    -- CP-element group 23: 	142 
    -- CP-element group 23: 	187 
    -- CP-element group 23: 	191 
    -- CP-element group 23: 	179 
    -- CP-element group 23: 	195 
    -- CP-element group 23: 	199 
    -- CP-element group 23: 	183 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/$entry
      -- CP-element group 23: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_6200_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	255 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	51 
    -- CP-element group 24: 	70 
    -- CP-element group 24: 	89 
    -- CP-element group 24: 	108 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/condition_evaluated
      -- 
    condition_evaluated_6318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(24), ack => do_while_stmt_2455_branch_req_0); -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(255) & convolve_CP_6200_elements(28) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(108);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	46 
    -- CP-element group 25: 	84 
    -- CP-element group 25: 	65 
    -- CP-element group 25: 	103 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	48 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	86 
    -- CP-element group 25: 	105 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/aggregated_phi_sample_req
      -- CP-element group 25: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_sample_start__ps
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(29) & convolve_CP_6200_elements(46) & convolve_CP_6200_elements(84) & convolve_CP_6200_elements(65) & convolve_CP_6200_elements(103) & convolve_CP_6200_elements(28);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	49 
    -- CP-element group 26: 	68 
    -- CP-element group 26: 	87 
    -- CP-element group 26: 	106 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	256 
    -- CP-element group 26: 	123 
    -- CP-element group 26: 	127 
    -- CP-element group 26: 	131 
    -- CP-element group 26: 	135 
    -- CP-element group 26: 	139 
    -- CP-element group 26: 	143 
    -- CP-element group 26: 	147 
    -- CP-element group 26: 	151 
    -- CP-element group 26: 	155 
    -- CP-element group 26: 	216 
    -- CP-element group 26: 	188 
    -- CP-element group 26: 	192 
    -- CP-element group 26: 	196 
    -- CP-element group 26: 	208 
    -- CP-element group 26: 	212 
    -- CP-element group 26: 	200 
    -- CP-element group 26: 	204 
    -- CP-element group 26: 	180 
    -- CP-element group 26: 	184 
    -- CP-element group 26: 	241 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	46 
    -- CP-element group 26: 	84 
    -- CP-element group 26: 	65 
    -- CP-element group 26: 	103 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/aggregated_phi_sample_ack
      -- CP-element group 26: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_sample_completed_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(31) & convolve_CP_6200_elements(49) & convolve_CP_6200_elements(68) & convolve_CP_6200_elements(87) & convolve_CP_6200_elements(106);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	47 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	85 
    -- CP-element group 27: 	104 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	50 
    -- CP-element group 27: 	69 
    -- CP-element group 27: 	88 
    -- CP-element group 27: 	107 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/aggregated_phi_update_req
      -- CP-element group 27: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_update_start__ps
      -- 
    convolve_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(30) & convolve_CP_6200_elements(47) & convolve_CP_6200_elements(66) & convolve_CP_6200_elements(85) & convolve_CP_6200_elements(104);
      gj_convolve_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	32 
    -- CP-element group 28: 	51 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	89 
    -- CP-element group 28: 	108 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(32) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(108);
      gj_convolve_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	125 
    -- CP-element group 29: 	129 
    -- CP-element group 29: 	133 
    -- CP-element group 29: 	137 
    -- CP-element group 29: 	141 
    -- CP-element group 29: 	145 
    -- CP-element group 29: 	149 
    -- CP-element group 29: 	153 
    -- CP-element group 29: 	157 
    -- CP-element group 29: 	214 
    -- CP-element group 29: 	218 
    -- CP-element group 29: 	186 
    -- CP-element group 29: 	190 
    -- CP-element group 29: 	194 
    -- CP-element group 29: 	198 
    -- CP-element group 29: 	206 
    -- CP-element group 29: 	210 
    -- CP-element group 29: 	202 
    -- CP-element group 29: 	182 
    -- CP-element group 29: 	243 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_sample_start_
      -- 
    convolve_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(26) & convolve_CP_6200_elements(125) & convolve_CP_6200_elements(129) & convolve_CP_6200_elements(133) & convolve_CP_6200_elements(137) & convolve_CP_6200_elements(141) & convolve_CP_6200_elements(145) & convolve_CP_6200_elements(149) & convolve_CP_6200_elements(153) & convolve_CP_6200_elements(157) & convolve_CP_6200_elements(214) & convolve_CP_6200_elements(218) & convolve_CP_6200_elements(186) & convolve_CP_6200_elements(190) & convolve_CP_6200_elements(194) & convolve_CP_6200_elements(198) & convolve_CP_6200_elements(206) & convolve_CP_6200_elements(210) & convolve_CP_6200_elements(202) & convolve_CP_6200_elements(182) & convolve_CP_6200_elements(243);
      gj_convolve_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	217 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	27 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_update_start_
      -- 
    convolve_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(32) & convolve_CP_6200_elements(217);
      gj_convolve_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_sample_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	28 
    -- CP-element group 32: 	215 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_update_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	21 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_loopback_trigger
      -- 
    convolve_CP_6200_elements(33) <= convolve_CP_6200_elements(21);
    -- CP-element group 34:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_loopback_sample_req
      -- CP-element group 34: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_loopback_sample_req_ps
      -- 
    phi_stmt_2457_loopback_sample_req_6333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2457_loopback_sample_req_6333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(34), ack => phi_stmt_2457_req_1); -- 
    -- Element group convolve_CP_6200_elements(34) is bound as output of CP function.
    -- CP-element group 35:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	22 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_entry_trigger
      -- 
    convolve_CP_6200_elements(35) <= convolve_CP_6200_elements(22);
    -- CP-element group 36:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_entry_sample_req
      -- CP-element group 36: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_entry_sample_req_ps
      -- 
    phi_stmt_2457_entry_sample_req_6336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2457_entry_sample_req_6336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(36), ack => phi_stmt_2457_req_0); -- 
    -- Element group convolve_CP_6200_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_phi_mux_ack
      -- CP-element group 37: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2457_phi_mux_ack_ps
      -- 
    phi_stmt_2457_phi_mux_ack_6339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2457_ack_0, ack => convolve_CP_6200_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_sample_completed_
      -- 
    -- Element group convolve_CP_6200_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_update_start_
      -- 
    -- Element group convolve_CP_6200_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_update_completed__ps
      -- 
    convolve_CP_6200_elements(40) <= convolve_CP_6200_elements(41);
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	40 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2461_update_completed_
      -- 
    -- Element group convolve_CP_6200_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => convolve_CP_6200_elements(39), ack => convolve_CP_6200_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_sample_start__ps
      -- CP-element group 42: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Sample/req
      -- 
    req_6360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(42), ack => nacc_2794_2462_buf_req_0); -- 
    -- Element group convolve_CP_6200_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_update_start__ps
      -- CP-element group 43: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_update_start_
      -- CP-element group 43: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Update/req
      -- 
    req_6365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(43), ack => nacc_2794_2462_buf_req_1); -- 
    -- Element group convolve_CP_6200_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_sample_completed__ps
      -- CP-element group 44: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Sample/ack
      -- 
    ack_6361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_2794_2462_buf_ack_0, ack => convolve_CP_6200_elements(44)); -- 
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_update_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_nacc_2462_Update/ack
      -- 
    ack_6366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_2794_2462_buf_ack_1, ack => convolve_CP_6200_elements(45)); -- 
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	26 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	25 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_sample_start_
      -- 
    convolve_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(26);
      gj_convolve_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	23 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	51 
    -- CP-element group 47: 	213 
    -- CP-element group 47: 	188 
    -- CP-element group 47: 	192 
    -- CP-element group 47: 	196 
    -- CP-element group 47: 	209 
    -- CP-element group 47: 	221 
    -- CP-element group 47: 	235 
    -- CP-element group 47: 	200 
    -- CP-element group 47: 	205 
    -- CP-element group 47: 	180 
    -- CP-element group 47: 	184 
    -- CP-element group 47: 	228 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	27 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_update_start_
      -- 
    convolve_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(213) & convolve_CP_6200_elements(188) & convolve_CP_6200_elements(192) & convolve_CP_6200_elements(196) & convolve_CP_6200_elements(209) & convolve_CP_6200_elements(221) & convolve_CP_6200_elements(235) & convolve_CP_6200_elements(200) & convolve_CP_6200_elements(205) & convolve_CP_6200_elements(180) & convolve_CP_6200_elements(184) & convolve_CP_6200_elements(228);
      gj_convolve_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	25 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_sample_start__ps
      -- 
    convolve_CP_6200_elements(48) <= convolve_CP_6200_elements(25);
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	26 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_sample_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	27 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_update_start__ps
      -- 
    convolve_CP_6200_elements(50) <= convolve_CP_6200_elements(27);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	24 
    -- CP-element group 51: 	28 
    -- CP-element group 51: 	219 
    -- CP-element group 51: 	188 
    -- CP-element group 51: 	192 
    -- CP-element group 51: 	196 
    -- CP-element group 51: 	207 
    -- CP-element group 51: 	211 
    -- CP-element group 51: 	233 
    -- CP-element group 51: 	200 
    -- CP-element group 51: 	203 
    -- CP-element group 51: 	180 
    -- CP-element group 51: 	184 
    -- CP-element group 51: 	226 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	47 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_update_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	21 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_loopback_trigger
      -- 
    convolve_CP_6200_elements(52) <= convolve_CP_6200_elements(21);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_loopback_sample_req
      -- CP-element group 53: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_loopback_sample_req_ps
      -- 
    phi_stmt_2463_loopback_sample_req_6377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2463_loopback_sample_req_6377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(53), ack => phi_stmt_2463_req_1); -- 
    -- Element group convolve_CP_6200_elements(53) is bound as output of CP function.
    -- CP-element group 54:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	22 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_entry_trigger
      -- 
    convolve_CP_6200_elements(54) <= convolve_CP_6200_elements(22);
    -- CP-element group 55:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_entry_sample_req
      -- CP-element group 55: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_entry_sample_req_ps
      -- 
    phi_stmt_2463_entry_sample_req_6380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2463_entry_sample_req_6380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(55), ack => phi_stmt_2463_req_0); -- 
    -- Element group convolve_CP_6200_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_phi_mux_ack
      -- CP-element group 56: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2463_phi_mux_ack_ps
      -- 
    phi_stmt_2463_phi_mux_ack_6383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2463_ack_0, ack => convolve_CP_6200_elements(56)); -- 
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_sample_start__ps
      -- CP-element group 57: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_sample_start_
      -- 
    -- Element group convolve_CP_6200_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_update_start_
      -- CP-element group 58: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_update_start__ps
      -- 
    -- Element group convolve_CP_6200_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_update_completed__ps
      -- 
    convolve_CP_6200_elements(59) <= convolve_CP_6200_elements(60);
    -- CP-element group 60:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	59 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2466_update_completed_
      -- 
    -- Element group convolve_CP_6200_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => convolve_CP_6200_elements(58), ack => convolve_CP_6200_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Sample/req
      -- CP-element group 61: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_sample_start__ps
      -- CP-element group 61: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_sample_start_
      -- 
    req_6404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(61), ack => n_row_2785_2467_buf_req_0); -- 
    -- Element group convolve_CP_6200_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_update_start__ps
      -- CP-element group 62: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Update/req
      -- CP-element group 62: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_update_start_
      -- 
    req_6409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(62), ack => n_row_2785_2467_buf_req_1); -- 
    -- Element group convolve_CP_6200_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_sample_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_sample_completed_
      -- 
    ack_6405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2785_2467_buf_ack_0, ack => convolve_CP_6200_elements(63)); -- 
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_update_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_row_2467_Update/$exit
      -- 
    ack_6410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2785_2467_buf_ack_1, ack => convolve_CP_6200_elements(64)); -- 
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	23 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	26 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	25 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_sample_start_
      -- 
    convolve_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(26);
      gj_convolve_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	23 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	70 
    -- CP-element group 66: 	123 
    -- CP-element group 66: 	127 
    -- CP-element group 66: 	131 
    -- CP-element group 66: 	135 
    -- CP-element group 66: 	139 
    -- CP-element group 66: 	143 
    -- CP-element group 66: 	148 
    -- CP-element group 66: 	152 
    -- CP-element group 66: 	156 
    -- CP-element group 66: 	160 
    -- CP-element group 66: 	213 
    -- CP-element group 66: 	167 
    -- CP-element group 66: 	188 
    -- CP-element group 66: 	192 
    -- CP-element group 66: 	174 
    -- CP-element group 66: 	196 
    -- CP-element group 66: 	209 
    -- CP-element group 66: 	221 
    -- CP-element group 66: 	235 
    -- CP-element group 66: 	200 
    -- CP-element group 66: 	205 
    -- CP-element group 66: 	180 
    -- CP-element group 66: 	184 
    -- CP-element group 66: 	228 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	27 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_update_start_
      -- 
    convolve_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 25) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1);
      constant place_markings: IntegerArray(0 to 25)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1);
      constant place_delays: IntegerArray(0 to 25) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 26); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(123) & convolve_CP_6200_elements(127) & convolve_CP_6200_elements(131) & convolve_CP_6200_elements(135) & convolve_CP_6200_elements(139) & convolve_CP_6200_elements(143) & convolve_CP_6200_elements(148) & convolve_CP_6200_elements(152) & convolve_CP_6200_elements(156) & convolve_CP_6200_elements(160) & convolve_CP_6200_elements(213) & convolve_CP_6200_elements(167) & convolve_CP_6200_elements(188) & convolve_CP_6200_elements(192) & convolve_CP_6200_elements(174) & convolve_CP_6200_elements(196) & convolve_CP_6200_elements(209) & convolve_CP_6200_elements(221) & convolve_CP_6200_elements(235) & convolve_CP_6200_elements(200) & convolve_CP_6200_elements(205) & convolve_CP_6200_elements(180) & convolve_CP_6200_elements(184) & convolve_CP_6200_elements(228);
      gj_convolve_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 26, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_sample_start__ps
      -- 
    convolve_CP_6200_elements(67) <= convolve_CP_6200_elements(25);
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	26 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_sample_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(68) is bound as output of CP function.
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	27 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_update_start__ps
      -- 
    convolve_CP_6200_elements(69) <= convolve_CP_6200_elements(27);
    -- CP-element group 70:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	24 
    -- CP-element group 70: 	28 
    -- CP-element group 70: 	123 
    -- CP-element group 70: 	127 
    -- CP-element group 70: 	131 
    -- CP-element group 70: 	135 
    -- CP-element group 70: 	139 
    -- CP-element group 70: 	143 
    -- CP-element group 70: 	146 
    -- CP-element group 70: 	150 
    -- CP-element group 70: 	154 
    -- CP-element group 70: 	158 
    -- CP-element group 70: 	219 
    -- CP-element group 70: 	165 
    -- CP-element group 70: 	188 
    -- CP-element group 70: 	192 
    -- CP-element group 70: 	196 
    -- CP-element group 70: 	172 
    -- CP-element group 70: 	207 
    -- CP-element group 70: 	211 
    -- CP-element group 70: 	233 
    -- CP-element group 70: 	200 
    -- CP-element group 70: 	203 
    -- CP-element group 70: 	180 
    -- CP-element group 70: 	184 
    -- CP-element group 70: 	226 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	66 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_update_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(70) is bound as output of CP function.
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	21 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_loopback_trigger
      -- 
    convolve_CP_6200_elements(71) <= convolve_CP_6200_elements(21);
    -- CP-element group 72:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_loopback_sample_req
      -- CP-element group 72: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_loopback_sample_req_ps
      -- 
    phi_stmt_2468_loopback_sample_req_6421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2468_loopback_sample_req_6421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(72), ack => phi_stmt_2468_req_1); -- 
    -- Element group convolve_CP_6200_elements(72) is bound as output of CP function.
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	22 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_entry_trigger
      -- 
    convolve_CP_6200_elements(73) <= convolve_CP_6200_elements(22);
    -- CP-element group 74:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_entry_sample_req
      -- CP-element group 74: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_entry_sample_req_ps
      -- 
    phi_stmt_2468_entry_sample_req_6424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2468_entry_sample_req_6424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(74), ack => phi_stmt_2468_req_0); -- 
    -- Element group convolve_CP_6200_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_phi_mux_ack
      -- CP-element group 75: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2468_phi_mux_ack_ps
      -- 
    phi_stmt_2468_phi_mux_ack_6427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2468_ack_0, ack => convolve_CP_6200_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_sample_start__ps
      -- CP-element group 76: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_sample_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_update_start__ps
      -- CP-element group 77: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_update_start_
      -- 
    -- Element group convolve_CP_6200_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_update_completed__ps
      -- 
    convolve_CP_6200_elements(78) <= convolve_CP_6200_elements(79);
    -- CP-element group 79:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	78 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2471_update_completed_
      -- 
    -- Element group convolve_CP_6200_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convolve_CP_6200_elements(77), ack => convolve_CP_6200_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_sample_start__ps
      -- CP-element group 80: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Sample/req
      -- 
    req_6448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(80), ack => n_col_2777_2472_buf_req_0); -- 
    -- Element group convolve_CP_6200_elements(80) is bound as output of CP function.
    -- CP-element group 81:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Update/req
      -- CP-element group 81: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_update_start__ps
      -- CP-element group 81: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_update_start_
      -- 
    req_6453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(81), ack => n_col_2777_2472_buf_req_1); -- 
    -- Element group convolve_CP_6200_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_sample_completed__ps
      -- CP-element group 82: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Sample/ack
      -- CP-element group 82: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_sample_completed_
      -- 
    ack_6449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2777_2472_buf_ack_0, ack => convolve_CP_6200_elements(82)); -- 
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Update/ack
      -- CP-element group 83: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_update_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_col_2472_Update/$exit
      -- 
    ack_6454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2777_2472_buf_ack_1, ack => convolve_CP_6200_elements(83)); -- 
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	23 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	26 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	25 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_sample_start_
      -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(26);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	23 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	89 
    -- CP-element group 85: 	123 
    -- CP-element group 85: 	127 
    -- CP-element group 85: 	131 
    -- CP-element group 85: 	135 
    -- CP-element group 85: 	139 
    -- CP-element group 85: 	143 
    -- CP-element group 85: 	148 
    -- CP-element group 85: 	152 
    -- CP-element group 85: 	156 
    -- CP-element group 85: 	160 
    -- CP-element group 85: 	167 
    -- CP-element group 85: 	174 
    -- CP-element group 85: 	242 
    -- CP-element group 85: 	246 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	27 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_update_start_
      -- 
    convolve_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(123) & convolve_CP_6200_elements(127) & convolve_CP_6200_elements(131) & convolve_CP_6200_elements(135) & convolve_CP_6200_elements(139) & convolve_CP_6200_elements(143) & convolve_CP_6200_elements(148) & convolve_CP_6200_elements(152) & convolve_CP_6200_elements(156) & convolve_CP_6200_elements(160) & convolve_CP_6200_elements(167) & convolve_CP_6200_elements(174) & convolve_CP_6200_elements(242) & convolve_CP_6200_elements(246);
      gj_convolve_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_sample_start__ps
      -- 
    convolve_CP_6200_elements(86) <= convolve_CP_6200_elements(25);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	26 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_sample_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(87) is bound as output of CP function.
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	27 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_update_start__ps
      -- 
    convolve_CP_6200_elements(88) <= convolve_CP_6200_elements(27);
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	24 
    -- CP-element group 89: 	28 
    -- CP-element group 89: 	123 
    -- CP-element group 89: 	127 
    -- CP-element group 89: 	131 
    -- CP-element group 89: 	135 
    -- CP-element group 89: 	139 
    -- CP-element group 89: 	143 
    -- CP-element group 89: 	146 
    -- CP-element group 89: 	150 
    -- CP-element group 89: 	154 
    -- CP-element group 89: 	158 
    -- CP-element group 89: 	165 
    -- CP-element group 89: 	172 
    -- CP-element group 89: 	240 
    -- CP-element group 89: 	244 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	85 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_update_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_update_completed_
      -- 
    -- Element group convolve_CP_6200_elements(89) is bound as output of CP function.
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	21 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_loopback_trigger
      -- 
    convolve_CP_6200_elements(90) <= convolve_CP_6200_elements(21);
    -- CP-element group 91:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_loopback_sample_req
      -- CP-element group 91: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_loopback_sample_req_ps
      -- 
    phi_stmt_2473_loopback_sample_req_6465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2473_loopback_sample_req_6465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(91), ack => phi_stmt_2473_req_1); -- 
    -- Element group convolve_CP_6200_elements(91) is bound as output of CP function.
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	22 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_entry_trigger
      -- 
    convolve_CP_6200_elements(92) <= convolve_CP_6200_elements(22);
    -- CP-element group 93:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_entry_sample_req
      -- CP-element group 93: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_entry_sample_req_ps
      -- 
    phi_stmt_2473_entry_sample_req_6468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2473_entry_sample_req_6468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(93), ack => phi_stmt_2473_req_0); -- 
    -- Element group convolve_CP_6200_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_phi_mux_ack
      -- CP-element group 94: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2473_phi_mux_ack_ps
      -- 
    phi_stmt_2473_phi_mux_ack_6471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2473_ack_0, ack => convolve_CP_6200_elements(94)); -- 
    -- CP-element group 95:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_sample_start__ps
      -- CP-element group 95: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_sample_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(95) is bound as output of CP function.
    -- CP-element group 96:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_update_start__ps
      -- CP-element group 96: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_update_start_
      -- 
    -- Element group convolve_CP_6200_elements(96) is bound as output of CP function.
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_update_completed__ps
      -- 
    convolve_CP_6200_elements(97) <= convolve_CP_6200_elements(98);
    -- CP-element group 98:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	97 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2477_update_completed_
      -- 
    -- Element group convolve_CP_6200_elements(98) is a control-delay.
    cp_element_98_delay: control_delay_element  generic map(name => " 98_delay", delay_value => 1)  port map(req => convolve_CP_6200_elements(96), ack => convolve_CP_6200_elements(98), clk => clk, reset =>reset);
    -- CP-element group 99:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (4) 
      -- CP-element group 99: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_sample_start__ps
      -- CP-element group 99: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Sample/req
      -- CP-element group 99: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_sample_start_
      -- 
    req_6492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(99), ack => n_num_2766_2478_buf_req_0); -- 
    -- Element group convolve_CP_6200_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_update_start__ps
      -- CP-element group 100: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Update/$entry
      -- 
    req_6497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(100), ack => n_num_2766_2478_buf_req_1); -- 
    -- Element group convolve_CP_6200_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_sample_completed__ps
      -- CP-element group 101: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Sample/ack
      -- 
    ack_6493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2766_2478_buf_ack_0, ack => convolve_CP_6200_elements(101)); -- 
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Update/ack
      -- CP-element group 102: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_num_2478_Update/$exit
      -- 
    ack_6498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2766_2478_buf_ack_1, ack => convolve_CP_6200_elements(102)); -- 
    -- CP-element group 103:  join  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	23 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	26 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	25 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_sample_start_
      -- 
    convolve_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(26);
      gj_convolve_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	23 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	108 
    -- CP-element group 104: 	242 
    -- CP-element group 104: 	246 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	27 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_update_start_
      -- 
    convolve_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(108) & convolve_CP_6200_elements(242) & convolve_CP_6200_elements(246);
      gj_convolve_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	25 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_sample_start__ps
      -- 
    convolve_CP_6200_elements(105) <= convolve_CP_6200_elements(25);
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	26 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_sample_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(106) is bound as output of CP function.
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	27 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_update_start__ps
      -- 
    convolve_CP_6200_elements(107) <= convolve_CP_6200_elements(27);
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	24 
    -- CP-element group 108: 	28 
    -- CP-element group 108: 	240 
    -- CP-element group 108: 	244 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	104 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_update_completed__ps
      -- 
    -- Element group convolve_CP_6200_elements(108) is bound as output of CP function.
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	21 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_loopback_trigger
      -- 
    convolve_CP_6200_elements(109) <= convolve_CP_6200_elements(21);
    -- CP-element group 110:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_loopback_sample_req_ps
      -- CP-element group 110: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_loopback_sample_req
      -- 
    phi_stmt_2479_loopback_sample_req_6509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2479_loopback_sample_req_6509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(110), ack => phi_stmt_2479_req_1); -- 
    -- Element group convolve_CP_6200_elements(110) is bound as output of CP function.
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	22 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_entry_trigger
      -- 
    convolve_CP_6200_elements(111) <= convolve_CP_6200_elements(22);
    -- CP-element group 112:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_entry_sample_req
      -- CP-element group 112: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_entry_sample_req_ps
      -- 
    phi_stmt_2479_entry_sample_req_6512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2479_entry_sample_req_6512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(112), ack => phi_stmt_2479_req_0); -- 
    -- Element group convolve_CP_6200_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_phi_mux_ack
      -- CP-element group 113: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/phi_stmt_2479_phi_mux_ack_ps
      -- 
    phi_stmt_2479_phi_mux_ack_6515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2479_ack_0, ack => convolve_CP_6200_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_sample_completed_
      -- 
    -- Element group convolve_CP_6200_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_update_start_
      -- 
    -- Element group convolve_CP_6200_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_update_completed__ps
      -- 
    convolve_CP_6200_elements(116) <= convolve_CP_6200_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2482_update_completed_
      -- 
    -- Element group convolve_CP_6200_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convolve_CP_6200_elements(115), ack => convolve_CP_6200_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Sample/req
      -- CP-element group 118: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_sample_start__ps
      -- 
    req_6536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(118), ack => n_chl_2755_2483_buf_req_0); -- 
    -- Element group convolve_CP_6200_elements(118) is bound as output of CP function.
    -- CP-element group 119:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_update_start_
      -- CP-element group 119: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_update_start__ps
      -- CP-element group 119: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Update/req
      -- 
    req_6541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(119), ack => n_chl_2755_2483_buf_req_1); -- 
    -- Element group convolve_CP_6200_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_sample_completed__ps
      -- 
    ack_6537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2755_2483_buf_ack_0, ack => convolve_CP_6200_elements(120)); -- 
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/R_n_chl_2483_Update/ack
      -- 
    ack_6542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2755_2483_buf_ack_1, ack => convolve_CP_6200_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	23 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	125 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Sample/rr
      -- 
    rr_6551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(122), ack => RPIPE_input_pipe1_2496_inst_req_0); -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(125);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	26 
    -- CP-element group 123: 	70 
    -- CP-element group 123: 	89 
    -- CP-element group 123: 	124 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	250 
    -- CP-element group 123: 	163 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	66 
    -- CP-element group 123: 	85 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_update_start_
      -- CP-element group 123: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Update/cr
      -- 
    cr_6556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(123), ack => RPIPE_input_pipe1_2496_inst_req_1); -- 
    convolve_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(124) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(163);
      gj_convolve_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Sample/ra
      -- 
    ra_6552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2496_inst_ack_0, ack => convolve_CP_6200_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	162 
    -- CP-element group 125: 	248 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	29 
    -- CP-element group 125: 	122 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe1_2496_Update/ca
      -- 
    ca_6557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2496_inst_ack_1, ack => convolve_CP_6200_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	23 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	129 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Sample/rr
      -- 
    rr_6565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(126), ack => RPIPE_input_pipe2_2500_inst_req_0); -- 
    convolve_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(129);
      gj_convolve_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	26 
    -- CP-element group 127: 	70 
    -- CP-element group 127: 	89 
    -- CP-element group 127: 	128 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	250 
    -- CP-element group 127: 	170 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	66 
    -- CP-element group 127: 	85 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_update_start_
      -- CP-element group 127: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Update/cr
      -- 
    cr_6570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(127), ack => RPIPE_input_pipe2_2500_inst_req_1); -- 
    convolve_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(128) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(170);
      gj_convolve_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	127 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Sample/ra
      -- 
    ra_6566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2500_inst_ack_0, ack => convolve_CP_6200_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	169 
    -- CP-element group 129: 	248 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	29 
    -- CP-element group 129: 	126 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe2_2500_Update/ca
      -- 
    ca_6571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2500_inst_ack_1, ack => convolve_CP_6200_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	23 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	133 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Sample/rr
      -- 
    rr_6579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(130), ack => RPIPE_input_pipe3_2504_inst_req_0); -- 
    convolve_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(133);
      gj_convolve_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	26 
    -- CP-element group 131: 	70 
    -- CP-element group 131: 	89 
    -- CP-element group 131: 	132 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	250 
    -- CP-element group 131: 	177 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	66 
    -- CP-element group 131: 	85 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_update_start_
      -- CP-element group 131: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Update/cr
      -- 
    cr_6584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(131), ack => RPIPE_input_pipe3_2504_inst_req_1); -- 
    convolve_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(132) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(177);
      gj_convolve_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	131 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Sample/ra
      -- 
    ra_6580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2504_inst_ack_0, ack => convolve_CP_6200_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	176 
    -- CP-element group 133: 	248 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	29 
    -- CP-element group 133: 	130 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_input_pipe3_2504_Update/ca
      -- 
    ca_6585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2504_inst_ack_1, ack => convolve_CP_6200_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	23 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	137 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Sample/rr
      -- 
    rr_6593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(134), ack => RPIPE_xxconvolvexxconv_ip1_2508_inst_req_0); -- 
    convolve_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(137);
      gj_convolve_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	26 
    -- CP-element group 135: 	70 
    -- CP-element group 135: 	89 
    -- CP-element group 135: 	136 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	250 
    -- CP-element group 135: 	163 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	66 
    -- CP-element group 135: 	85 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_update_start_
      -- CP-element group 135: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Update/cr
      -- 
    cr_6598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(135), ack => RPIPE_xxconvolvexxconv_ip1_2508_inst_req_1); -- 
    convolve_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(136) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(163);
      gj_convolve_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Sample/ra
      -- 
    ra_6594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2508_inst_ack_0, ack => convolve_CP_6200_elements(136)); -- 
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	162 
    -- CP-element group 137: 	248 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	29 
    -- CP-element group 137: 	134 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip1_2508_Update/ca
      -- 
    ca_6599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2508_inst_ack_1, ack => convolve_CP_6200_elements(137)); -- 
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	23 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	141 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Sample/rr
      -- 
    rr_6607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(138), ack => RPIPE_xxconvolvexxconv_ip2_2512_inst_req_0); -- 
    convolve_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(141);
      gj_convolve_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	26 
    -- CP-element group 139: 	70 
    -- CP-element group 139: 	89 
    -- CP-element group 139: 	140 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	250 
    -- CP-element group 139: 	170 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	66 
    -- CP-element group 139: 	85 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_update_start_
      -- CP-element group 139: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Update/cr
      -- 
    cr_6612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(139), ack => RPIPE_xxconvolvexxconv_ip2_2512_inst_req_1); -- 
    convolve_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(140) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(170);
      gj_convolve_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	139 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Sample/ra
      -- 
    ra_6608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2512_inst_ack_0, ack => convolve_CP_6200_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	169 
    -- CP-element group 141: 	248 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	29 
    -- CP-element group 141: 	138 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip2_2512_Update/ca
      -- 
    ca_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2512_inst_ack_1, ack => convolve_CP_6200_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	23 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	145 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Sample/rr
      -- 
    rr_6621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(142), ack => RPIPE_xxconvolvexxconv_ip3_2516_inst_req_0); -- 
    convolve_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(145);
      gj_convolve_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	26 
    -- CP-element group 143: 	70 
    -- CP-element group 143: 	89 
    -- CP-element group 143: 	144 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	250 
    -- CP-element group 143: 	177 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	66 
    -- CP-element group 143: 	85 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_update_start_
      -- CP-element group 143: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Update/cr
      -- 
    cr_6626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(143), ack => RPIPE_xxconvolvexxconv_ip3_2516_inst_req_1); -- 
    convolve_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(144) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(177);
      gj_convolve_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	143 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Sample/ra
      -- 
    ra_6622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2516_inst_ack_0, ack => convolve_CP_6200_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	176 
    -- CP-element group 145: 	248 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	29 
    -- CP-element group 145: 	142 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_ip3_2516_Update/ca
      -- 
    ca_6627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2516_inst_ack_1, ack => convolve_CP_6200_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	70 
    -- CP-element group 146: 	89 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Sample/req
      -- 
    req_6635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(146), ack => W_read_ip_2474_delayed_1_0_2518_inst_req_0); -- 
    convolve_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(148);
      gj_convolve_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	26 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	250 
    -- CP-element group 147: 	149 
    -- CP-element group 147: 	163 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_update_start_
      -- CP-element group 147: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Update/req
      -- 
    req_6640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(147), ack => W_read_ip_2474_delayed_1_0_2518_inst_req_1); -- 
    convolve_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(149) & convolve_CP_6200_elements(163);
      gj_convolve_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	66 
    -- CP-element group 148: 	85 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Sample/ack
      -- 
    ack_6636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2474_delayed_1_0_2518_inst_ack_0, ack => convolve_CP_6200_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	162 
    -- CP-element group 149: 	248 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	29 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2520_Update/ack
      -- 
    ack_6641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2474_delayed_1_0_2518_inst_ack_1, ack => convolve_CP_6200_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	70 
    -- CP-element group 150: 	89 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Sample/req
      -- 
    req_6649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(150), ack => W_read_ip_2480_delayed_1_0_2527_inst_req_0); -- 
    convolve_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(152);
      gj_convolve_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	26 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	250 
    -- CP-element group 151: 	153 
    -- CP-element group 151: 	170 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_update_start_
      -- CP-element group 151: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Update/req
      -- 
    req_6654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(151), ack => W_read_ip_2480_delayed_1_0_2527_inst_req_1); -- 
    convolve_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(153) & convolve_CP_6200_elements(170);
      gj_convolve_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	66 
    -- CP-element group 152: 	85 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Sample/ack
      -- 
    ack_6650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2480_delayed_1_0_2527_inst_ack_0, ack => convolve_CP_6200_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	169 
    -- CP-element group 153: 	248 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	29 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2529_Update/ack
      -- 
    ack_6655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2480_delayed_1_0_2527_inst_ack_1, ack => convolve_CP_6200_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	70 
    -- CP-element group 154: 	89 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Sample/req
      -- 
    req_6663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(154), ack => W_read_ip_2486_delayed_1_0_2536_inst_req_0); -- 
    convolve_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(156);
      gj_convolve_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	26 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	250 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	177 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_update_start_
      -- CP-element group 155: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Update/req
      -- 
    req_6668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(155), ack => W_read_ip_2486_delayed_1_0_2536_inst_req_1); -- 
    convolve_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(157) & convolve_CP_6200_elements(177);
      gj_convolve_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	66 
    -- CP-element group 156: 	85 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Sample/ack
      -- 
    ack_6664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2486_delayed_1_0_2536_inst_ack_0, ack => convolve_CP_6200_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	176 
    -- CP-element group 157: 	248 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	29 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2538_Update/ack
      -- 
    ack_6669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2486_delayed_1_0_2536_inst_ack_1, ack => convolve_CP_6200_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	70 
    -- CP-element group 158: 	89 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Sample/req
      -- 
    req_6677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(158), ack => W_write_input_2500_delayed_1_0_2554_inst_req_0); -- 
    convolve_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(160);
      gj_convolve_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: 	163 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_update_start_
      -- CP-element group 159: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Update/req
      -- 
    req_6682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(159), ack => W_write_input_2500_delayed_1_0_2554_inst_req_1); -- 
    convolve_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(161) & convolve_CP_6200_elements(163);
      gj_convolve_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	66 
    -- CP-element group 160: 	85 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Sample/ack
      -- 
    ack_6678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2500_delayed_1_0_2554_inst_ack_0, ack => convolve_CP_6200_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2556_Update/ack
      -- 
    ack_6683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2500_delayed_1_0_2554_inst_ack_1, ack => convolve_CP_6200_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	125 
    -- CP-element group 162: 	137 
    -- CP-element group 162: 	149 
    -- CP-element group 162: 	161 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Sample/req
      -- 
    req_6691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(162), ack => WPIPE_xxconvolvexxconv_ip1_2558_inst_req_0); -- 
    convolve_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(125) & convolve_CP_6200_elements(137) & convolve_CP_6200_elements(149) & convolve_CP_6200_elements(161) & convolve_CP_6200_elements(164);
      gj_convolve_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	123 
    -- CP-element group 163: 	135 
    -- CP-element group 163: 	147 
    -- CP-element group 163: 	159 
    -- CP-element group 163:  members (6) 
      -- CP-element group 163: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_update_start_
      -- CP-element group 163: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Sample/ack
      -- CP-element group 163: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Update/req
      -- 
    ack_6692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2558_inst_ack_0, ack => convolve_CP_6200_elements(163)); -- 
    req_6696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(163), ack => WPIPE_xxconvolvexxconv_ip1_2558_inst_req_1); -- 
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	256 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip1_2558_Update/ack
      -- 
    ack_6697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2558_inst_ack_1, ack => convolve_CP_6200_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	70 
    -- CP-element group 165: 	89 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Sample/req
      -- 
    req_6705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(165), ack => W_write_input_2504_delayed_1_0_2561_inst_req_0); -- 
    convolve_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(167);
      gj_convolve_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: 	170 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_update_start_
      -- CP-element group 166: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Update/req
      -- 
    req_6710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(166), ack => W_write_input_2504_delayed_1_0_2561_inst_req_1); -- 
    convolve_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(168) & convolve_CP_6200_elements(170);
      gj_convolve_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	66 
    -- CP-element group 167: 	85 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Sample/ack
      -- 
    ack_6706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2504_delayed_1_0_2561_inst_ack_0, ack => convolve_CP_6200_elements(167)); -- 
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2563_Update/ack
      -- 
    ack_6711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2504_delayed_1_0_2561_inst_ack_1, ack => convolve_CP_6200_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	129 
    -- CP-element group 169: 	141 
    -- CP-element group 169: 	153 
    -- CP-element group 169: 	168 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Sample/req
      -- 
    req_6719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(169), ack => WPIPE_xxconvolvexxconv_ip2_2565_inst_req_0); -- 
    convolve_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(129) & convolve_CP_6200_elements(141) & convolve_CP_6200_elements(153) & convolve_CP_6200_elements(168) & convolve_CP_6200_elements(171);
      gj_convolve_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	127 
    -- CP-element group 170: 	139 
    -- CP-element group 170: 	151 
    -- CP-element group 170: 	166 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_update_start_
      -- CP-element group 170: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Sample/ack
      -- CP-element group 170: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Update/req
      -- 
    ack_6720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2565_inst_ack_0, ack => convolve_CP_6200_elements(170)); -- 
    req_6724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(170), ack => WPIPE_xxconvolvexxconv_ip2_2565_inst_req_1); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	256 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip2_2565_Update/ack
      -- 
    ack_6725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2565_inst_ack_1, ack => convolve_CP_6200_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	70 
    -- CP-element group 172: 	89 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Sample/req
      -- 
    req_6733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(172), ack => W_write_input_2508_delayed_1_0_2568_inst_req_0); -- 
    convolve_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(70) & convolve_CP_6200_elements(89) & convolve_CP_6200_elements(174);
      gj_convolve_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	177 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_update_start_
      -- CP-element group 173: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Update/req
      -- 
    req_6738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(173), ack => W_write_input_2508_delayed_1_0_2568_inst_req_1); -- 
    convolve_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(175) & convolve_CP_6200_elements(177);
      gj_convolve_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	66 
    -- CP-element group 174: 	85 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Sample/ack
      -- 
    ack_6734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2508_delayed_1_0_2568_inst_ack_0, ack => convolve_CP_6200_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2570_Update/ack
      -- 
    ack_6739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2508_delayed_1_0_2568_inst_ack_1, ack => convolve_CP_6200_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	133 
    -- CP-element group 176: 	145 
    -- CP-element group 176: 	157 
    -- CP-element group 176: 	175 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Sample/req
      -- 
    req_6747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(176), ack => WPIPE_xxconvolvexxconv_ip3_2572_inst_req_0); -- 
    convolve_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(133) & convolve_CP_6200_elements(145) & convolve_CP_6200_elements(157) & convolve_CP_6200_elements(175) & convolve_CP_6200_elements(178);
      gj_convolve_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	131 
    -- CP-element group 177: 	143 
    -- CP-element group 177: 	155 
    -- CP-element group 177: 	173 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_update_start_
      -- CP-element group 177: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Sample/ack
      -- CP-element group 177: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Update/req
      -- 
    ack_6748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2572_inst_ack_0, ack => convolve_CP_6200_elements(177)); -- 
    req_6752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(177), ack => WPIPE_xxconvolvexxconv_ip3_2572_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	256 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_ip3_2572_Update/ack
      -- 
    ack_6753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2572_inst_ack_1, ack => convolve_CP_6200_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	23 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	182 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Sample/rr
      -- 
    rr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(179), ack => RPIPE_kernel_pipe1_2598_inst_req_0); -- 
    convolve_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(182);
      gj_convolve_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	26 
    -- CP-element group 180: 	51 
    -- CP-element group 180: 	70 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	250 
    -- CP-element group 180: 	224 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	47 
    -- CP-element group 180: 	66 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_update_start_
      -- CP-element group 180: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Update/cr
      -- 
    cr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(180), ack => RPIPE_kernel_pipe1_2598_inst_req_1); -- 
    convolve_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(181) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(224);
      gj_convolve_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	180 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Sample/ra
      -- 
    ra_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2598_inst_ack_0, ack => convolve_CP_6200_elements(181)); -- 
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	223 
    -- CP-element group 182: 	248 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	29 
    -- CP-element group 182: 	179 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe1_2598_Update/ca
      -- 
    ca_6767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2598_inst_ack_1, ack => convolve_CP_6200_elements(182)); -- 
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	23 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	186 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Sample/rr
      -- 
    rr_6775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(183), ack => RPIPE_kernel_pipe2_2602_inst_req_0); -- 
    convolve_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(186);
      gj_convolve_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	26 
    -- CP-element group 184: 	51 
    -- CP-element group 184: 	70 
    -- CP-element group 184: 	185 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	250 
    -- CP-element group 184: 	231 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	47 
    -- CP-element group 184: 	66 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_update_start_
      -- CP-element group 184: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Update/cr
      -- 
    cr_6780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(184), ack => RPIPE_kernel_pipe2_2602_inst_req_1); -- 
    convolve_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(185) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(231);
      gj_convolve_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	184 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Sample/ra
      -- 
    ra_6776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2602_inst_ack_0, ack => convolve_CP_6200_elements(185)); -- 
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	230 
    -- CP-element group 186: 	248 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	29 
    -- CP-element group 186: 	183 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe2_2602_Update/ca
      -- 
    ca_6781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2602_inst_ack_1, ack => convolve_CP_6200_elements(186)); -- 
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	23 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	190 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Sample/rr
      -- 
    rr_6789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(187), ack => RPIPE_kernel_pipe3_2606_inst_req_0); -- 
    convolve_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(190);
      gj_convolve_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	26 
    -- CP-element group 188: 	51 
    -- CP-element group 188: 	70 
    -- CP-element group 188: 	189 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	250 
    -- CP-element group 188: 	238 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	47 
    -- CP-element group 188: 	66 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_update_start_
      -- CP-element group 188: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Update/cr
      -- 
    cr_6794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(188), ack => RPIPE_kernel_pipe3_2606_inst_req_1); -- 
    convolve_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(189) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(238);
      gj_convolve_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	188 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Sample/ra
      -- 
    ra_6790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2606_inst_ack_0, ack => convolve_CP_6200_elements(189)); -- 
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	237 
    -- CP-element group 190: 	248 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	29 
    -- CP-element group 190: 	187 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_kernel_pipe3_2606_Update/ca
      -- 
    ca_6795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2606_inst_ack_1, ack => convolve_CP_6200_elements(190)); -- 
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	23 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	194 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Sample/rr
      -- 
    rr_6803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(191), ack => RPIPE_xxconvolvexxconv_k1_2610_inst_req_0); -- 
    convolve_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(194);
      gj_convolve_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	26 
    -- CP-element group 192: 	51 
    -- CP-element group 192: 	70 
    -- CP-element group 192: 	193 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	250 
    -- CP-element group 192: 	224 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	47 
    -- CP-element group 192: 	66 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_update_start_
      -- CP-element group 192: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Update/$entry
      -- CP-element group 192: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Update/cr
      -- 
    cr_6808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(192), ack => RPIPE_xxconvolvexxconv_k1_2610_inst_req_1); -- 
    convolve_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(193) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(224);
      gj_convolve_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	192 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Sample/ra
      -- 
    ra_6804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2610_inst_ack_0, ack => convolve_CP_6200_elements(193)); -- 
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	223 
    -- CP-element group 194: 	248 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	29 
    -- CP-element group 194: 	191 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k1_2610_Update/ca
      -- 
    ca_6809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2610_inst_ack_1, ack => convolve_CP_6200_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	23 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	198 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Sample/rr
      -- 
    rr_6817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(195), ack => RPIPE_xxconvolvexxconv_k2_2614_inst_req_0); -- 
    convolve_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(198);
      gj_convolve_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	26 
    -- CP-element group 196: 	51 
    -- CP-element group 196: 	70 
    -- CP-element group 196: 	197 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	250 
    -- CP-element group 196: 	231 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	47 
    -- CP-element group 196: 	66 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_update_start_
      -- CP-element group 196: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Update/$entry
      -- CP-element group 196: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Update/cr
      -- 
    cr_6822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(196), ack => RPIPE_xxconvolvexxconv_k2_2614_inst_req_1); -- 
    convolve_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(197) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(231);
      gj_convolve_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	196 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Sample/ra
      -- 
    ra_6818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2614_inst_ack_0, ack => convolve_CP_6200_elements(197)); -- 
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	230 
    -- CP-element group 198: 	248 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	29 
    -- CP-element group 198: 	195 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k2_2614_Update/ca
      -- 
    ca_6823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2614_inst_ack_1, ack => convolve_CP_6200_elements(198)); -- 
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	23 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	202 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Sample/rr
      -- 
    rr_6831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(199), ack => RPIPE_xxconvolvexxconv_k3_2618_inst_req_0); -- 
    convolve_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(23) & convolve_CP_6200_elements(202);
      gj_convolve_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	26 
    -- CP-element group 200: 	51 
    -- CP-element group 200: 	70 
    -- CP-element group 200: 	201 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	250 
    -- CP-element group 200: 	238 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	47 
    -- CP-element group 200: 	66 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_update_start_
      -- CP-element group 200: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Update/cr
      -- 
    cr_6836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(200), ack => RPIPE_xxconvolvexxconv_k3_2618_inst_req_1); -- 
    convolve_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(201) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(238);
      gj_convolve_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	200 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Sample/ra
      -- 
    ra_6832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2618_inst_ack_0, ack => convolve_CP_6200_elements(201)); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	237 
    -- CP-element group 202: 	248 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	29 
    -- CP-element group 202: 	199 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/RPIPE_xxconvolvexxconv_k3_2618_Update/ca
      -- 
    ca_6837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2618_inst_ack_1, ack => convolve_CP_6200_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	51 
    -- CP-element group 203: 	70 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Sample/req
      -- 
    req_6845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(203), ack => W_read_k_2558_delayed_1_0_2620_inst_req_0); -- 
    convolve_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(205);
      gj_convolve_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	26 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	250 
    -- CP-element group 204: 	206 
    -- CP-element group 204: 	224 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_update_start_
      -- CP-element group 204: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Update/req
      -- 
    req_6850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(204), ack => W_read_k_2558_delayed_1_0_2620_inst_req_1); -- 
    convolve_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(206) & convolve_CP_6200_elements(224);
      gj_convolve_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	47 
    -- CP-element group 205: 	66 
    -- CP-element group 205: 	203 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Sample/ack
      -- 
    ack_6846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2558_delayed_1_0_2620_inst_ack_0, ack => convolve_CP_6200_elements(205)); -- 
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	223 
    -- CP-element group 206: 	248 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	29 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2622_Update/ack
      -- 
    ack_6851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2558_delayed_1_0_2620_inst_ack_1, ack => convolve_CP_6200_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	51 
    -- CP-element group 207: 	70 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Sample/req
      -- 
    req_6859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(207), ack => W_read_k_2564_delayed_1_0_2629_inst_req_0); -- 
    convolve_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(209);
      gj_convolve_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	26 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	250 
    -- CP-element group 208: 	210 
    -- CP-element group 208: 	231 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_update_start_
      -- CP-element group 208: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Update/req
      -- 
    req_6864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(208), ack => W_read_k_2564_delayed_1_0_2629_inst_req_1); -- 
    convolve_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(210) & convolve_CP_6200_elements(231);
      gj_convolve_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	47 
    -- CP-element group 209: 	66 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Sample/ack
      -- 
    ack_6860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2564_delayed_1_0_2629_inst_ack_0, ack => convolve_CP_6200_elements(209)); -- 
    -- CP-element group 210:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	230 
    -- CP-element group 210: 	248 
    -- CP-element group 210: marked-successors 
    -- CP-element group 210: 	29 
    -- CP-element group 210: 	208 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2631_Update/ack
      -- 
    ack_6865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2564_delayed_1_0_2629_inst_ack_1, ack => convolve_CP_6200_elements(210)); -- 
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	51 
    -- CP-element group 211: 	70 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Sample/req
      -- 
    req_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(211), ack => W_read_k_2570_delayed_1_0_2638_inst_req_0); -- 
    convolve_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(213);
      gj_convolve_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	26 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	250 
    -- CP-element group 212: 	214 
    -- CP-element group 212: 	238 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_update_start_
      -- CP-element group 212: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Update/req
      -- 
    req_6878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(212), ack => W_read_k_2570_delayed_1_0_2638_inst_req_1); -- 
    convolve_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(214) & convolve_CP_6200_elements(238);
      gj_convolve_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	47 
    -- CP-element group 213: 	66 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Sample/ack
      -- 
    ack_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2570_delayed_1_0_2638_inst_ack_0, ack => convolve_CP_6200_elements(213)); -- 
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	237 
    -- CP-element group 214: 	248 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	29 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2640_Update/ack
      -- 
    ack_6879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2570_delayed_1_0_2638_inst_ack_1, ack => convolve_CP_6200_elements(214)); -- 
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	32 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	217 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Sample/req
      -- 
    req_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(215), ack => W_acc_2606_delayed_1_0_2677_inst_req_0); -- 
    convolve_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(32) & convolve_CP_6200_elements(217);
      gj_convolve_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	26 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	250 
    -- CP-element group 216: 	218 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_update_start_
      -- CP-element group 216: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Update/req
      -- 
    req_6892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(216), ack => W_acc_2606_delayed_1_0_2677_inst_req_1); -- 
    convolve_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(250) & convolve_CP_6200_elements(218);
      gj_convolve_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: marked-successors 
    -- CP-element group 217: 	30 
    -- CP-element group 217: 	215 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Sample/ack
      -- 
    ack_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_2606_delayed_1_0_2677_inst_ack_0, ack => convolve_CP_6200_elements(217)); -- 
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	248 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	29 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2679_Update/ack
      -- 
    ack_6893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_2606_delayed_1_0_2677_inst_ack_1, ack => convolve_CP_6200_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	51 
    -- CP-element group 219: 	70 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Sample/req
      -- 
    req_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(219), ack => W_store_kernel_2652_delayed_1_0_2727_inst_req_0); -- 
    convolve_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(221);
      gj_convolve_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: 	224 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_update_start_
      -- CP-element group 220: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Update/req
      -- 
    req_6906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(220), ack => W_store_kernel_2652_delayed_1_0_2727_inst_req_1); -- 
    convolve_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(222) & convolve_CP_6200_elements(224);
      gj_convolve_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: marked-successors 
    -- CP-element group 221: 	47 
    -- CP-element group 221: 	66 
    -- CP-element group 221: 	219 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Sample/ack
      -- 
    ack_6902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2652_delayed_1_0_2727_inst_ack_0, ack => convolve_CP_6200_elements(221)); -- 
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2729_Update/ack
      -- 
    ack_6907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2652_delayed_1_0_2727_inst_ack_1, ack => convolve_CP_6200_elements(222)); -- 
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	194 
    -- CP-element group 223: 	206 
    -- CP-element group 223: 	222 
    -- CP-element group 223: 	182 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	225 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Sample/req
      -- 
    req_6915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(223), ack => WPIPE_xxconvolvexxconv_k1_2731_inst_req_0); -- 
    convolve_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(194) & convolve_CP_6200_elements(206) & convolve_CP_6200_elements(222) & convolve_CP_6200_elements(182) & convolve_CP_6200_elements(225);
      gj_convolve_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	192 
    -- CP-element group 224: 	220 
    -- CP-element group 224: 	204 
    -- CP-element group 224: 	180 
    -- CP-element group 224:  members (6) 
      -- CP-element group 224: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_update_start_
      -- CP-element group 224: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Sample/ack
      -- CP-element group 224: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Update/req
      -- 
    ack_6916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2731_inst_ack_0, ack => convolve_CP_6200_elements(224)); -- 
    req_6920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(224), ack => WPIPE_xxconvolvexxconv_k1_2731_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	256 
    -- CP-element group 225: marked-successors 
    -- CP-element group 225: 	223 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k1_2731_Update/ack
      -- 
    ack_6921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2731_inst_ack_1, ack => convolve_CP_6200_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	51 
    -- CP-element group 226: 	70 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Sample/req
      -- 
    req_6929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(226), ack => W_store_kernel_2656_delayed_1_0_2734_inst_req_0); -- 
    convolve_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(228);
      gj_convolve_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	231 
    -- CP-element group 227: 	229 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Update/req
      -- CP-element group 227: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_update_start_
      -- 
    req_6934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(227), ack => W_store_kernel_2656_delayed_1_0_2734_inst_req_1); -- 
    convolve_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(231) & convolve_CP_6200_elements(229);
      gj_convolve_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	47 
    -- CP-element group 228: 	66 
    -- CP-element group 228: 	226 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Sample/ack
      -- CP-element group 228: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_sample_completed_
      -- 
    ack_6930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2656_delayed_1_0_2734_inst_ack_0, ack => convolve_CP_6200_elements(228)); -- 
    -- CP-element group 229:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229: marked-successors 
    -- CP-element group 229: 	227 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Update/ack
      -- CP-element group 229: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2736_update_completed_
      -- 
    ack_6935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2656_delayed_1_0_2734_inst_ack_1, ack => convolve_CP_6200_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	186 
    -- CP-element group 230: 	198 
    -- CP-element group 230: 	210 
    -- CP-element group 230: 	229 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Sample/req
      -- 
    req_6943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(230), ack => WPIPE_xxconvolvexxconv_k2_2738_inst_req_0); -- 
    convolve_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(186) & convolve_CP_6200_elements(198) & convolve_CP_6200_elements(210) & convolve_CP_6200_elements(229) & convolve_CP_6200_elements(232);
      gj_convolve_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	196 
    -- CP-element group 231: 	208 
    -- CP-element group 231: 	184 
    -- CP-element group 231: 	227 
    -- CP-element group 231:  members (6) 
      -- CP-element group 231: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Update/req
      -- CP-element group 231: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_update_start_
      -- CP-element group 231: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Sample/ack
      -- 
    ack_6944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2738_inst_ack_0, ack => convolve_CP_6200_elements(231)); -- 
    req_6948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(231), ack => WPIPE_xxconvolvexxconv_k2_2738_inst_req_1); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	256 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Update/ack
      -- CP-element group 232: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k2_2738_Update/$exit
      -- 
    ack_6949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2738_inst_ack_1, ack => convolve_CP_6200_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	51 
    -- CP-element group 233: 	70 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Sample/req
      -- 
    req_6957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(233), ack => W_store_kernel_2660_delayed_1_0_2741_inst_req_0); -- 
    convolve_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(51) & convolve_CP_6200_elements(70) & convolve_CP_6200_elements(235);
      gj_convolve_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: 	238 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_update_start_
      -- CP-element group 234: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Update/req
      -- 
    req_6962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(234), ack => W_store_kernel_2660_delayed_1_0_2741_inst_req_1); -- 
    convolve_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(236) & convolve_CP_6200_elements(238);
      gj_convolve_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	47 
    -- CP-element group 235: 	66 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Sample/$exit
      -- 
    ack_6958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2660_delayed_1_0_2741_inst_ack_0, ack => convolve_CP_6200_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2743_Update/ack
      -- 
    ack_6963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2660_delayed_1_0_2741_inst_ack_1, ack => convolve_CP_6200_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	214 
    -- CP-element group 237: 	190 
    -- CP-element group 237: 	236 
    -- CP-element group 237: 	202 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Sample/req
      -- CP-element group 237: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Sample/$entry
      -- 
    req_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(237), ack => WPIPE_xxconvolvexxconv_k3_2745_inst_req_0); -- 
    convolve_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(214) & convolve_CP_6200_elements(190) & convolve_CP_6200_elements(236) & convolve_CP_6200_elements(202) & convolve_CP_6200_elements(239);
      gj_convolve_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	188 
    -- CP-element group 238: 	212 
    -- CP-element group 238: 	234 
    -- CP-element group 238: 	200 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Update/req
      -- CP-element group 238: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Sample/ack
      -- CP-element group 238: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_update_start_
      -- CP-element group 238: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_sample_completed_
      -- 
    ack_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2745_inst_ack_0, ack => convolve_CP_6200_elements(238)); -- 
    req_6976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(238), ack => WPIPE_xxconvolvexxconv_k3_2745_inst_req_1); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	256 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Update/ack
      -- CP-element group 239: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_xxconvolvexxconv_k3_2745_update_completed_
      -- 
    ack_6977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2745_inst_ack_1, ack => convolve_CP_6200_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	89 
    -- CP-element group 240: 	108 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	242 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Sample/req
      -- 
    req_6985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(240), ack => W_num_done_2703_delayed_1_0_2786_inst_req_0); -- 
    convolve_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(89) & convolve_CP_6200_elements(108) & convolve_CP_6200_elements(242);
      gj_convolve_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	26 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_update_start_
      -- CP-element group 241: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Update/req
      -- 
    req_6990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(241), ack => W_num_done_2703_delayed_1_0_2786_inst_req_1); -- 
    convolve_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(26) & convolve_CP_6200_elements(243);
      gj_convolve_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: marked-successors 
    -- CP-element group 242: 	85 
    -- CP-element group 242: 	104 
    -- CP-element group 242: 	240 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Sample/ack
      -- CP-element group 242: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_sample_completed_
      -- 
    ack_6986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2703_delayed_1_0_2786_inst_ack_0, ack => convolve_CP_6200_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	256 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	29 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_Update/ack
      -- CP-element group 243: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2788_update_completed_
      -- 
    ack_6991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2703_delayed_1_0_2786_inst_ack_1, ack => convolve_CP_6200_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	89 
    -- CP-element group 244: 	108 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Sample/$entry
      -- 
    req_6999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(244), ack => W_num_done_2708_delayed_1_0_2795_inst_req_0); -- 
    convolve_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(89) & convolve_CP_6200_elements(108) & convolve_CP_6200_elements(246);
      gj_convolve_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	250 
    -- CP-element group 245: 	253 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Update/req
      -- CP-element group 245: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_update_start_
      -- 
    req_7004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(245), ack => W_num_done_2708_delayed_1_0_2795_inst_req_1); -- 
    convolve_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(250) & convolve_CP_6200_elements(253) & convolve_CP_6200_elements(247);
      gj_convolve_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	85 
    -- CP-element group 246: 	104 
    -- CP-element group 246: 	244 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Sample/ack
      -- CP-element group 246: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_sample_completed_
      -- 
    ack_7000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2708_delayed_1_0_2795_inst_ack_0, ack => convolve_CP_6200_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	252 
    -- CP-element group 247: 	248 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Update/ack
      -- CP-element group 247: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/assign_stmt_2797_update_completed_
      -- 
    ack_7005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2708_delayed_1_0_2795_inst_ack_1, ack => convolve_CP_6200_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	125 
    -- CP-element group 248: 	129 
    -- CP-element group 248: 	133 
    -- CP-element group 248: 	137 
    -- CP-element group 248: 	141 
    -- CP-element group 248: 	145 
    -- CP-element group 248: 	149 
    -- CP-element group 248: 	153 
    -- CP-element group 248: 	157 
    -- CP-element group 248: 	214 
    -- CP-element group 248: 	218 
    -- CP-element group 248: 	186 
    -- CP-element group 248: 	190 
    -- CP-element group 248: 	194 
    -- CP-element group 248: 	198 
    -- CP-element group 248: 	206 
    -- CP-element group 248: 	210 
    -- CP-element group 248: 	202 
    -- CP-element group 248: 	182 
    -- CP-element group 248: 	247 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Sample/rr
      -- 
    rr_7013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(248), ack => type_cast_2801_inst_req_0); -- 
    convolve_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(125) & convolve_CP_6200_elements(129) & convolve_CP_6200_elements(133) & convolve_CP_6200_elements(137) & convolve_CP_6200_elements(141) & convolve_CP_6200_elements(145) & convolve_CP_6200_elements(149) & convolve_CP_6200_elements(153) & convolve_CP_6200_elements(157) & convolve_CP_6200_elements(214) & convolve_CP_6200_elements(218) & convolve_CP_6200_elements(186) & convolve_CP_6200_elements(190) & convolve_CP_6200_elements(194) & convolve_CP_6200_elements(198) & convolve_CP_6200_elements(206) & convolve_CP_6200_elements(210) & convolve_CP_6200_elements(202) & convolve_CP_6200_elements(182) & convolve_CP_6200_elements(247) & convolve_CP_6200_elements(250);
      gj_convolve_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	253 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_update_start_
      -- 
    cr_7018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(249), ack => type_cast_2801_inst_req_1); -- 
    convolve_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(251) & convolve_CP_6200_elements(253);
      gj_convolve_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	123 
    -- CP-element group 250: 	127 
    -- CP-element group 250: 	131 
    -- CP-element group 250: 	135 
    -- CP-element group 250: 	139 
    -- CP-element group 250: 	143 
    -- CP-element group 250: 	147 
    -- CP-element group 250: 	151 
    -- CP-element group 250: 	155 
    -- CP-element group 250: 	216 
    -- CP-element group 250: 	188 
    -- CP-element group 250: 	192 
    -- CP-element group 250: 	196 
    -- CP-element group 250: 	208 
    -- CP-element group 250: 	212 
    -- CP-element group 250: 	200 
    -- CP-element group 250: 	204 
    -- CP-element group 250: 	180 
    -- CP-element group 250: 	184 
    -- CP-element group 250: 	245 
    -- CP-element group 250: 	248 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Sample/ra
      -- CP-element group 250: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Sample/$exit
      -- 
    ra_7014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2801_inst_ack_0, ack => convolve_CP_6200_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/type_cast_2801_Update/ca
      -- 
    ca_7019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2801_inst_ack_1, ack => convolve_CP_6200_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: 	247 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_sample_start_
      -- 
    req_7027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(252), ack => WPIPE_output_pipe_2799_inst_req_0); -- 
    convolve_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(251) & convolve_CP_6200_elements(247) & convolve_CP_6200_elements(254);
      gj_convolve_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253: marked-successors 
    -- CP-element group 253: 	245 
    -- CP-element group 253: 	249 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_update_start_
      -- CP-element group 253: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Update/req
      -- CP-element group 253: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_sample_completed_
      -- 
    ack_7028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2799_inst_ack_0, ack => convolve_CP_6200_elements(253)); -- 
    req_7032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(253), ack => WPIPE_output_pipe_2799_inst_req_1); -- 
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/WPIPE_output_pipe_2799_Update/$exit
      -- 
    ack_7033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2799_inst_ack_1, ack => convolve_CP_6200_elements(254)); -- 
    -- CP-element group 255:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	23 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	24 
    -- CP-element group 255:  members (1) 
      -- CP-element group 255: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_6200_elements(255) is a control-delay.
    cp_element_255_delay: control_delay_element  generic map(name => " 255_delay", delay_value => 1)  port map(req => convolve_CP_6200_elements(23), ack => convolve_CP_6200_elements(255), clk => clk, reset =>reset);
    -- CP-element group 256:  join  transition  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	26 
    -- CP-element group 256: 	164 
    -- CP-element group 256: 	178 
    -- CP-element group 256: 	171 
    -- CP-element group 256: 	232 
    -- CP-element group 256: 	225 
    -- CP-element group 256: 	239 
    -- CP-element group 256: 	243 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	20 
    -- CP-element group 256:  members (1) 
      -- CP-element group 256: 	 branch_block_stmt_2438/do_while_stmt_2455/do_while_stmt_2455_loop_body/$exit
      -- 
    convolve_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolve_CP_6200_elements(254) & convolve_CP_6200_elements(26) & convolve_CP_6200_elements(164) & convolve_CP_6200_elements(178) & convolve_CP_6200_elements(171) & convolve_CP_6200_elements(232) & convolve_CP_6200_elements(225) & convolve_CP_6200_elements(239) & convolve_CP_6200_elements(243);
      gj_convolve_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6200_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	19 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (2) 
      -- CP-element group 257: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_exit/ack
      -- CP-element group 257: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_exit/$exit
      -- 
    ack_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2455_branch_ack_0, ack => convolve_CP_6200_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	19 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_taken/$exit
      -- CP-element group 258: 	 branch_block_stmt_2438/do_while_stmt_2455/loop_taken/ack
      -- 
    ack_7042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2455_branch_ack_1, ack => convolve_CP_6200_elements(258)); -- 
    -- CP-element group 259:  transition  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	17 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	2 
    -- CP-element group 259:  members (1) 
      -- CP-element group 259: 	 branch_block_stmt_2438/do_while_stmt_2455/$exit
      -- 
    convolve_CP_6200_elements(259) <= convolve_CP_6200_elements(17);
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	2 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_update_start_
      -- CP-element group 260: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Update/req
      -- CP-element group 260: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Sample/ack
      -- 
    ack_7055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_2806_inst_ack_0, ack => convolve_CP_6200_elements(260)); -- 
    req_7059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(260), ack => WPIPE_input_done_pipe_2806_inst_req_1); -- 
    -- CP-element group 261:  transition  place  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (8) 
      -- CP-element group 261: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Update/ack
      -- CP-element group 261: 	 branch_block_stmt_2438/loopback_PhiReq/$entry
      -- CP-element group 261: 	 branch_block_stmt_2438/loopback_PhiReq/$exit
      -- CP-element group 261: 	 branch_block_stmt_2438/assign_stmt_2808/$exit
      -- CP-element group 261: 	 branch_block_stmt_2438/assign_stmt_2808__exit__
      -- CP-element group 261: 	 branch_block_stmt_2438/loopback
      -- CP-element group 261: 	 branch_block_stmt_2438/assign_stmt_2808/WPIPE_input_done_pipe_2806_Update/$exit
      -- 
    ack_7060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_2806_inst_ack_1, ack => convolve_CP_6200_elements(261)); -- 
    -- CP-element group 262:  merge  fork  transition  place  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: 	0 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	10 
    -- CP-element group 262: 	11 
    -- CP-element group 262: 	14 
    -- CP-element group 262: 	3 
    -- CP-element group 262: 	6 
    -- CP-element group 262:  members (22) 
      -- CP-element group 262: 	 branch_block_stmt_2438/merge_stmt_2439_PhiReqMerge
      -- CP-element group 262: 	 branch_block_stmt_2438/merge_stmt_2439_PhiAck/dummy
      -- CP-element group 262: 	 branch_block_stmt_2438/merge_stmt_2439_PhiAck/$entry
      -- CP-element group 262: 	 branch_block_stmt_2438/merge_stmt_2439_PhiAck/$exit
      -- CP-element group 262: 	 branch_block_stmt_2438/merge_stmt_2439__exit__
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454__entry__
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/$entry
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_update_start_
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_num_out_pipe_2441_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2443_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_update_start_
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2448_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_update_start_
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/RPIPE_size_pipe_2451_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_2438/assign_stmt_2444_to_assign_stmt_2454/SUB_u16_u16_2453_Update/cr
      -- 
    rr_6231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(262), ack => RPIPE_num_out_pipe_2441_inst_req_0); -- 
    cr_6246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(262), ack => SUB_u16_u16_2443_inst_req_1); -- 
    cr_6274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(262), ack => SUB_u16_u16_2448_inst_req_1); -- 
    rr_6287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(262), ack => RPIPE_size_pipe_2451_inst_req_0); -- 
    cr_6302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6200_elements(262), ack => SUB_u16_u16_2453_inst_req_1); -- 
    convolve_CP_6200_elements(262) <= OrReduce(convolve_CP_6200_elements(261) & convolve_CP_6200_elements(0));
    convolve_do_while_stmt_2455_terminator_7043: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_2455_terminator_7043", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_6200_elements(20),loop_continue => convolve_CP_6200_elements(258),loop_terminate => convolve_CP_6200_elements(257),loop_back => convolve_CP_6200_elements(18),loop_exit => convolve_CP_6200_elements(17),clk => clk, reset => reset); -- 
    phi_stmt_2457_phi_seq_6367_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6200_elements(35);
      convolve_CP_6200_elements(38)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6200_elements(38);
      convolve_CP_6200_elements(39)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6200_elements(40);
      convolve_CP_6200_elements(36) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6200_elements(33);
      convolve_CP_6200_elements(42)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6200_elements(44);
      convolve_CP_6200_elements(43)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6200_elements(45);
      convolve_CP_6200_elements(34) <= phi_mux_reqs(1);
      phi_stmt_2457_phi_seq_6367 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2457_phi_seq_6367") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6200_elements(25), 
          phi_sample_ack => convolve_CP_6200_elements(31), 
          phi_update_req => convolve_CP_6200_elements(27), 
          phi_update_ack => convolve_CP_6200_elements(32), 
          phi_mux_ack => convolve_CP_6200_elements(37), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2463_phi_seq_6411_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6200_elements(54);
      convolve_CP_6200_elements(57)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6200_elements(57);
      convolve_CP_6200_elements(58)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6200_elements(59);
      convolve_CP_6200_elements(55) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6200_elements(52);
      convolve_CP_6200_elements(61)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6200_elements(63);
      convolve_CP_6200_elements(62)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6200_elements(64);
      convolve_CP_6200_elements(53) <= phi_mux_reqs(1);
      phi_stmt_2463_phi_seq_6411 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2463_phi_seq_6411") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6200_elements(48), 
          phi_sample_ack => convolve_CP_6200_elements(49), 
          phi_update_req => convolve_CP_6200_elements(50), 
          phi_update_ack => convolve_CP_6200_elements(51), 
          phi_mux_ack => convolve_CP_6200_elements(56), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2468_phi_seq_6455_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6200_elements(73);
      convolve_CP_6200_elements(76)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6200_elements(76);
      convolve_CP_6200_elements(77)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6200_elements(78);
      convolve_CP_6200_elements(74) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6200_elements(71);
      convolve_CP_6200_elements(80)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6200_elements(82);
      convolve_CP_6200_elements(81)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6200_elements(83);
      convolve_CP_6200_elements(72) <= phi_mux_reqs(1);
      phi_stmt_2468_phi_seq_6455 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2468_phi_seq_6455") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6200_elements(67), 
          phi_sample_ack => convolve_CP_6200_elements(68), 
          phi_update_req => convolve_CP_6200_elements(69), 
          phi_update_ack => convolve_CP_6200_elements(70), 
          phi_mux_ack => convolve_CP_6200_elements(75), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2473_phi_seq_6499_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6200_elements(92);
      convolve_CP_6200_elements(95)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6200_elements(95);
      convolve_CP_6200_elements(96)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6200_elements(97);
      convolve_CP_6200_elements(93) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6200_elements(90);
      convolve_CP_6200_elements(99)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6200_elements(101);
      convolve_CP_6200_elements(100)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6200_elements(102);
      convolve_CP_6200_elements(91) <= phi_mux_reqs(1);
      phi_stmt_2473_phi_seq_6499 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2473_phi_seq_6499") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6200_elements(86), 
          phi_sample_ack => convolve_CP_6200_elements(87), 
          phi_update_req => convolve_CP_6200_elements(88), 
          phi_update_ack => convolve_CP_6200_elements(89), 
          phi_mux_ack => convolve_CP_6200_elements(94), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2479_phi_seq_6543_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6200_elements(111);
      convolve_CP_6200_elements(114)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6200_elements(114);
      convolve_CP_6200_elements(115)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6200_elements(116);
      convolve_CP_6200_elements(112) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6200_elements(109);
      convolve_CP_6200_elements(118)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6200_elements(120);
      convolve_CP_6200_elements(119)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6200_elements(121);
      convolve_CP_6200_elements(110) <= phi_mux_reqs(1);
      phi_stmt_2479_phi_seq_6543 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2479_phi_seq_6543") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6200_elements(105), 
          phi_sample_ack => convolve_CP_6200_elements(106), 
          phi_update_req => convolve_CP_6200_elements(107), 
          phi_update_ack => convolve_CP_6200_elements(108), 
          phi_mux_ack => convolve_CP_6200_elements(113), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6319_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_6200_elements(21);
        preds(1)  <= convolve_CP_6200_elements(22);
        entry_tmerge_6319 : transition_merge -- 
          generic map(name => " entry_tmerge_6319")
          port map (preds => preds, symbol_out => convolve_CP_6200_elements(23));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_i16_i16_2683_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_2686_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2753_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2773_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2782_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_2762_wire : std_logic_vector(1 downto 0);
    signal AND_u1_u1_2719_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2488_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2590_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2593_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2491_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2697_wire : std_logic_vector(0 downto 0);
    signal MUL_i16_i16_2662_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2668_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2674_wire : std_logic_vector(15 downto 0);
    signal MUX_2763_wire : std_logic_vector(1 downto 0);
    signal MUX_2774_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_2805_wire : std_logic_vector(0 downto 0);
    signal RPIPE_num_out_pipe_2441_wire : std_logic_vector(15 downto 0);
    signal RPIPE_num_out_pipe_2446_wire : std_logic_vector(15 downto 0);
    signal RPIPE_size_pipe_2451_wire : std_logic_vector(15 downto 0);
    signal UGT_u2_u1_2551_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_2548_wire : std_logic_vector(0 downto 0);
    signal acc_2457 : std_logic_vector(15 downto 0);
    signal acc_2606_delayed_1_0_2679 : std_logic_vector(15 downto 0);
    signal acc_val_2688 : std_logic_vector(15 downto 0);
    signal all_done_flag_2726 : std_logic_vector(0 downto 0);
    signal chl_2479 : std_logic_vector(15 downto 0);
    signal chl_done_2693 : std_logic_vector(0 downto 0);
    signal col_2468 : std_logic_vector(15 downto 0);
    signal col_done_2705 : std_logic_vector(0 downto 0);
    signal iread1_2526 : std_logic_vector(15 downto 0);
    signal iread2_2535 : std_logic_vector(15 downto 0);
    signal iread3_2544 : std_logic_vector(15 downto 0);
    signal ival1_2578 : std_logic_vector(15 downto 0);
    signal ival2_2582 : std_logic_vector(15 downto 0);
    signal ival3_2586 : std_logic_vector(15 downto 0);
    signal konst_2442_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2447_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2452_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2487_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2490_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2550_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2589_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2592_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2696_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2750_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2752_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2759_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2761_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2770_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2772_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2781_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2791_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2807_wire_constant : std_logic_vector(7 downto 0);
    signal kread1_2628 : std_logic_vector(15 downto 0);
    signal kread2_2637 : std_logic_vector(15 downto 0);
    signal kread3_2646 : std_logic_vector(15 downto 0);
    signal kval1_2650 : std_logic_vector(15 downto 0);
    signal kval2_2654 : std_logic_vector(15 downto 0);
    signal kval3_2658 : std_logic_vector(15 downto 0);
    signal mul_val1_2664 : std_logic_vector(15 downto 0);
    signal mul_val2_2670 : std_logic_vector(15 downto 0);
    signal mul_val3_2676 : std_logic_vector(15 downto 0);
    signal n_chl_2755 : std_logic_vector(15 downto 0);
    signal n_chl_2755_2483_buffered : std_logic_vector(15 downto 0);
    signal n_col_2777 : std_logic_vector(15 downto 0);
    signal n_col_2777_2472_buffered : std_logic_vector(15 downto 0);
    signal n_num_2766 : std_logic_vector(1 downto 0);
    signal n_num_2766_2478_buffered : std_logic_vector(1 downto 0);
    signal n_row_2785 : std_logic_vector(15 downto 0);
    signal n_row_2785_2467_buffered : std_logic_vector(15 downto 0);
    signal nacc_2794 : std_logic_vector(15 downto 0);
    signal nacc_2794_2462_buffered : std_logic_vector(15 downto 0);
    signal num_2473 : std_logic_vector(1 downto 0);
    signal num_chl_2454 : std_logic_vector(15 downto 0);
    signal num_col_2449 : std_logic_vector(15 downto 0);
    signal num_done_2700 : std_logic_vector(0 downto 0);
    signal num_done_2703_delayed_1_0_2788 : std_logic_vector(0 downto 0);
    signal num_done_2708_delayed_1_0_2797 : std_logic_vector(0 downto 0);
    signal num_row_2444 : std_logic_vector(15 downto 0);
    signal out_done_flag_2715 : std_logic_vector(0 downto 0);
    signal read_ip_2474_delayed_1_0_2520 : std_logic_vector(0 downto 0);
    signal read_ip_2480_delayed_1_0_2529 : std_logic_vector(0 downto 0);
    signal read_ip_2486_delayed_1_0_2538 : std_logic_vector(0 downto 0);
    signal read_ip_2493 : std_logic_vector(0 downto 0);
    signal read_k_2558_delayed_1_0_2622 : std_logic_vector(0 downto 0);
    signal read_k_2564_delayed_1_0_2631 : std_logic_vector(0 downto 0);
    signal read_k_2570_delayed_1_0_2640 : std_logic_vector(0 downto 0);
    signal read_k_2595 : std_logic_vector(0 downto 0);
    signal row_2463 : std_logic_vector(15 downto 0);
    signal row_done_2710 : std_logic_vector(0 downto 0);
    signal store_kernel_2652_delayed_1_0_2729 : std_logic_vector(0 downto 0);
    signal store_kernel_2656_delayed_1_0_2736 : std_logic_vector(0 downto 0);
    signal store_kernel_2660_delayed_1_0_2743 : std_logic_vector(0 downto 0);
    signal store_kernel_2721 : std_logic_vector(0 downto 0);
    signal temp1_1_2509 : std_logic_vector(15 downto 0);
    signal temp1_2_2513 : std_logic_vector(15 downto 0);
    signal temp1_3_2517 : std_logic_vector(15 downto 0);
    signal temp2_1_2497 : std_logic_vector(15 downto 0);
    signal temp2_2_2501 : std_logic_vector(15 downto 0);
    signal temp2_3_2505 : std_logic_vector(15 downto 0);
    signal tempk1_1_2599 : std_logic_vector(15 downto 0);
    signal tempk1_2_2603 : std_logic_vector(15 downto 0);
    signal tempk1_3_2607 : std_logic_vector(15 downto 0);
    signal tempk2_1_2611 : std_logic_vector(15 downto 0);
    signal tempk2_2_2615 : std_logic_vector(15 downto 0);
    signal tempk2_3_2619 : std_logic_vector(15 downto 0);
    signal type_cast_2461_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2466_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2471_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2477_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_2482_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2801_wire : std_logic_vector(15 downto 0);
    signal write_input_2500_delayed_1_0_2556 : std_logic_vector(0 downto 0);
    signal write_input_2504_delayed_1_0_2563 : std_logic_vector(0 downto 0);
    signal write_input_2508_delayed_1_0_2570 : std_logic_vector(0 downto 0);
    signal write_input_2553 : std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_2442_wire_constant <= "0000000000000001";
    konst_2447_wire_constant <= "0000000000000001";
    konst_2452_wire_constant <= "0000000000000001";
    konst_2487_wire_constant <= "0000000000000000";
    konst_2490_wire_constant <= "10";
    konst_2550_wire_constant <= "00";
    konst_2589_wire_constant <= "0000000000000000";
    konst_2592_wire_constant <= "0000000000000000";
    konst_2696_wire_constant <= "10";
    konst_2750_wire_constant <= "0000000000000000";
    konst_2752_wire_constant <= "0000000000000001";
    konst_2759_wire_constant <= "00";
    konst_2761_wire_constant <= "01";
    konst_2770_wire_constant <= "0000000000000000";
    konst_2772_wire_constant <= "0000000000000001";
    konst_2781_wire_constant <= "0000000000000001";
    konst_2791_wire_constant <= "0000000000000000";
    konst_2807_wire_constant <= "00000001";
    type_cast_2461_wire_constant <= "0000000000000000";
    type_cast_2466_wire_constant <= "0000000000000000";
    type_cast_2471_wire_constant <= "0000000000000000";
    type_cast_2477_wire_constant <= "00";
    type_cast_2482_wire_constant <= "0000000000000000";
    phi_stmt_2457: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2461_wire_constant & nacc_2794_2462_buffered;
      req <= phi_stmt_2457_req_0 & phi_stmt_2457_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2457",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2457_ack_0,
          idata => idata,
          odata => acc_2457,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2457
    phi_stmt_2463: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2466_wire_constant & n_row_2785_2467_buffered;
      req <= phi_stmt_2463_req_0 & phi_stmt_2463_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2463",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2463_ack_0,
          idata => idata,
          odata => row_2463,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2463
    phi_stmt_2468: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2471_wire_constant & n_col_2777_2472_buffered;
      req <= phi_stmt_2468_req_0 & phi_stmt_2468_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2468",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2468_ack_0,
          idata => idata,
          odata => col_2468,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2468
    phi_stmt_2473: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2477_wire_constant & n_num_2766_2478_buffered;
      req <= phi_stmt_2473_req_0 & phi_stmt_2473_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2473",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2473_ack_0,
          idata => idata,
          odata => num_2473,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2473
    phi_stmt_2479: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2482_wire_constant & n_chl_2755_2483_buffered;
      req <= phi_stmt_2479_req_0 & phi_stmt_2479_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2479",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2479_ack_0,
          idata => idata,
          odata => chl_2479,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2479
    -- flow-through select operator MUX_2525_inst
    iread1_2526 <= temp2_1_2497 when (read_ip_2474_delayed_1_0_2520(0) /=  '0') else temp1_1_2509;
    -- flow-through select operator MUX_2534_inst
    iread2_2535 <= temp2_2_2501 when (read_ip_2480_delayed_1_0_2529(0) /=  '0') else temp1_2_2513;
    -- flow-through select operator MUX_2543_inst
    iread3_2544 <= temp2_3_2505 when (read_ip_2486_delayed_1_0_2538(0) /=  '0') else temp1_3_2517;
    -- flow-through select operator MUX_2627_inst
    kread1_2628 <= tempk1_1_2599 when (read_k_2558_delayed_1_0_2622(0) /=  '0') else tempk2_1_2611;
    -- flow-through select operator MUX_2636_inst
    kread2_2637 <= tempk1_2_2603 when (read_k_2564_delayed_1_0_2631(0) /=  '0') else tempk2_2_2615;
    -- flow-through select operator MUX_2645_inst
    kread3_2646 <= tempk1_3_2607 when (read_k_2570_delayed_1_0_2640(0) /=  '0') else tempk2_3_2619;
    -- flow-through select operator MUX_2754_inst
    n_chl_2755 <= konst_2750_wire_constant when (chl_done_2693(0) /=  '0') else ADD_u16_u16_2753_wire;
    -- flow-through select operator MUX_2763_inst
    MUX_2763_wire <= konst_2759_wire_constant when (num_done_2700(0) /=  '0') else ADD_u2_u2_2762_wire;
    -- flow-through select operator MUX_2765_inst
    n_num_2766 <= MUX_2763_wire when (chl_done_2693(0) /=  '0') else num_2473;
    -- flow-through select operator MUX_2774_inst
    MUX_2774_wire <= konst_2770_wire_constant when (col_done_2705(0) /=  '0') else ADD_u16_u16_2773_wire;
    -- flow-through select operator MUX_2776_inst
    n_col_2777 <= MUX_2774_wire when (num_done_2700(0) /=  '0') else col_2468;
    -- flow-through select operator MUX_2784_inst
    n_row_2785 <= ADD_u16_u16_2782_wire when (row_done_2710(0) /=  '0') else row_2463;
    -- flow-through select operator MUX_2793_inst
    nacc_2794 <= konst_2791_wire_constant when (num_done_2703_delayed_1_0_2788(0) /=  '0') else acc_val_2688;
    W_acc_2606_delayed_1_0_2677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc_2606_delayed_1_0_2677_inst_req_0;
      W_acc_2606_delayed_1_0_2677_inst_ack_0<= wack(0);
      rreq(0) <= W_acc_2606_delayed_1_0_2677_inst_req_1;
      W_acc_2606_delayed_1_0_2677_inst_ack_1<= rack(0);
      W_acc_2606_delayed_1_0_2677_inst : InterlockBuffer generic map ( -- 
        name => "W_acc_2606_delayed_1_0_2677_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_2457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc_2606_delayed_1_0_2679,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2703_delayed_1_0_2786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2703_delayed_1_0_2786_inst_req_0;
      W_num_done_2703_delayed_1_0_2786_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2703_delayed_1_0_2786_inst_req_1;
      W_num_done_2703_delayed_1_0_2786_inst_ack_1<= rack(0);
      W_num_done_2703_delayed_1_0_2786_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2703_delayed_1_0_2786_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2700,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2703_delayed_1_0_2788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2708_delayed_1_0_2795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2708_delayed_1_0_2795_inst_req_0;
      W_num_done_2708_delayed_1_0_2795_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2708_delayed_1_0_2795_inst_req_1;
      W_num_done_2708_delayed_1_0_2795_inst_ack_1<= rack(0);
      W_num_done_2708_delayed_1_0_2795_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2708_delayed_1_0_2795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2700,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2708_delayed_1_0_2797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2474_delayed_1_0_2518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2474_delayed_1_0_2518_inst_req_0;
      W_read_ip_2474_delayed_1_0_2518_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2474_delayed_1_0_2518_inst_req_1;
      W_read_ip_2474_delayed_1_0_2518_inst_ack_1<= rack(0);
      W_read_ip_2474_delayed_1_0_2518_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2474_delayed_1_0_2518_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2493,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2474_delayed_1_0_2520,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2480_delayed_1_0_2527_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2480_delayed_1_0_2527_inst_req_0;
      W_read_ip_2480_delayed_1_0_2527_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2480_delayed_1_0_2527_inst_req_1;
      W_read_ip_2480_delayed_1_0_2527_inst_ack_1<= rack(0);
      W_read_ip_2480_delayed_1_0_2527_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2480_delayed_1_0_2527_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2493,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2480_delayed_1_0_2529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2486_delayed_1_0_2536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2486_delayed_1_0_2536_inst_req_0;
      W_read_ip_2486_delayed_1_0_2536_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2486_delayed_1_0_2536_inst_req_1;
      W_read_ip_2486_delayed_1_0_2536_inst_ack_1<= rack(0);
      W_read_ip_2486_delayed_1_0_2536_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2486_delayed_1_0_2536_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2493,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2486_delayed_1_0_2538,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2558_delayed_1_0_2620_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2558_delayed_1_0_2620_inst_req_0;
      W_read_k_2558_delayed_1_0_2620_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2558_delayed_1_0_2620_inst_req_1;
      W_read_k_2558_delayed_1_0_2620_inst_ack_1<= rack(0);
      W_read_k_2558_delayed_1_0_2620_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2558_delayed_1_0_2620_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2558_delayed_1_0_2622,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2564_delayed_1_0_2629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2564_delayed_1_0_2629_inst_req_0;
      W_read_k_2564_delayed_1_0_2629_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2564_delayed_1_0_2629_inst_req_1;
      W_read_k_2564_delayed_1_0_2629_inst_ack_1<= rack(0);
      W_read_k_2564_delayed_1_0_2629_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2564_delayed_1_0_2629_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2564_delayed_1_0_2631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2570_delayed_1_0_2638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2570_delayed_1_0_2638_inst_req_0;
      W_read_k_2570_delayed_1_0_2638_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2570_delayed_1_0_2638_inst_req_1;
      W_read_k_2570_delayed_1_0_2638_inst_ack_1<= rack(0);
      W_read_k_2570_delayed_1_0_2638_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2570_delayed_1_0_2638_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2570_delayed_1_0_2640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2652_delayed_1_0_2727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2652_delayed_1_0_2727_inst_req_0;
      W_store_kernel_2652_delayed_1_0_2727_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2652_delayed_1_0_2727_inst_req_1;
      W_store_kernel_2652_delayed_1_0_2727_inst_ack_1<= rack(0);
      W_store_kernel_2652_delayed_1_0_2727_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2652_delayed_1_0_2727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2652_delayed_1_0_2729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2656_delayed_1_0_2734_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2656_delayed_1_0_2734_inst_req_0;
      W_store_kernel_2656_delayed_1_0_2734_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2656_delayed_1_0_2734_inst_req_1;
      W_store_kernel_2656_delayed_1_0_2734_inst_ack_1<= rack(0);
      W_store_kernel_2656_delayed_1_0_2734_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2656_delayed_1_0_2734_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2656_delayed_1_0_2736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2660_delayed_1_0_2741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2660_delayed_1_0_2741_inst_req_0;
      W_store_kernel_2660_delayed_1_0_2741_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2660_delayed_1_0_2741_inst_req_1;
      W_store_kernel_2660_delayed_1_0_2741_inst_ack_1<= rack(0);
      W_store_kernel_2660_delayed_1_0_2741_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2660_delayed_1_0_2741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2660_delayed_1_0_2743,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2500_delayed_1_0_2554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2500_delayed_1_0_2554_inst_req_0;
      W_write_input_2500_delayed_1_0_2554_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2500_delayed_1_0_2554_inst_req_1;
      W_write_input_2500_delayed_1_0_2554_inst_ack_1<= rack(0);
      W_write_input_2500_delayed_1_0_2554_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2500_delayed_1_0_2554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2500_delayed_1_0_2556,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2504_delayed_1_0_2561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2504_delayed_1_0_2561_inst_req_0;
      W_write_input_2504_delayed_1_0_2561_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2504_delayed_1_0_2561_inst_req_1;
      W_write_input_2504_delayed_1_0_2561_inst_ack_1<= rack(0);
      W_write_input_2504_delayed_1_0_2561_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2504_delayed_1_0_2561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2504_delayed_1_0_2563,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2508_delayed_1_0_2568_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2508_delayed_1_0_2568_inst_req_0;
      W_write_input_2508_delayed_1_0_2568_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2508_delayed_1_0_2568_inst_req_1;
      W_write_input_2508_delayed_1_0_2568_inst_ack_1<= rack(0);
      W_write_input_2508_delayed_1_0_2568_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2508_delayed_1_0_2568_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2508_delayed_1_0_2570,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_2755_2483_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_2755_2483_buf_req_0;
      n_chl_2755_2483_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_2755_2483_buf_req_1;
      n_chl_2755_2483_buf_ack_1<= rack(0);
      n_chl_2755_2483_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_2755_2483_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_2755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_2755_2483_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_2777_2472_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_2777_2472_buf_req_0;
      n_col_2777_2472_buf_ack_0<= wack(0);
      rreq(0) <= n_col_2777_2472_buf_req_1;
      n_col_2777_2472_buf_ack_1<= rack(0);
      n_col_2777_2472_buf : InterlockBuffer generic map ( -- 
        name => "n_col_2777_2472_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_2777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_2777_2472_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_num_2766_2478_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_num_2766_2478_buf_req_0;
      n_num_2766_2478_buf_ack_0<= wack(0);
      rreq(0) <= n_num_2766_2478_buf_req_1;
      n_num_2766_2478_buf_ack_1<= rack(0);
      n_num_2766_2478_buf : InterlockBuffer generic map ( -- 
        name => "n_num_2766_2478_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_num_2766,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_num_2766_2478_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_2785_2467_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_2785_2467_buf_req_0;
      n_row_2785_2467_buf_ack_0<= wack(0);
      rreq(0) <= n_row_2785_2467_buf_req_1;
      n_row_2785_2467_buf_ack_1<= rack(0);
      n_row_2785_2467_buf : InterlockBuffer generic map ( -- 
        name => "n_row_2785_2467_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_2785,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_2785_2467_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_2794_2462_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_2794_2462_buf_req_0;
      nacc_2794_2462_buf_ack_0<= wack(0);
      rreq(0) <= nacc_2794_2462_buf_req_1;
      nacc_2794_2462_buf_ack_1<= rack(0);
      nacc_2794_2462_buf : InterlockBuffer generic map ( -- 
        name => "nacc_2794_2462_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_2794,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_2794_2462_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2577_inst
    process(iread1_2526) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread1_2526(15 downto 0);
      ival1_2578 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2581_inst
    process(iread2_2535) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread2_2535(15 downto 0);
      ival2_2582 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2585_inst
    process(iread3_2544) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread3_2544(15 downto 0);
      ival3_2586 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2649_inst
    process(kread1_2628) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread1_2628(15 downto 0);
      kval1_2650 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2653_inst
    process(kread2_2637) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread2_2637(15 downto 0);
      kval2_2654 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2657_inst
    process(kread3_2646) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread3_2646(15 downto 0);
      kval3_2658 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2663_inst
    process(MUL_i16_i16_2662_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2662_wire(15 downto 0);
      mul_val1_2664 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2669_inst
    process(MUL_i16_i16_2668_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2668_wire(15 downto 0);
      mul_val2_2670 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2675_inst
    process(MUL_i16_i16_2674_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2674_wire(15 downto 0);
      mul_val3_2676 <= tmp_var; -- 
    end process;
    type_cast_2801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_2801_inst_req_0;
      type_cast_2801_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_2801_inst_req_1;
      type_cast_2801_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  num_done_2708_delayed_1_0_2797(0);
      type_cast_2801_inst_gI: SplitGuardInterface generic map(name => "type_cast_2801_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_2801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_2688,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2801_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_2455_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2805_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2455_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2455_branch_req_0,
          ack0 => do_while_stmt_2455_branch_ack_0,
          ack1 => do_while_stmt_2455_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_2683_inst
    process(acc_2606_delayed_1_0_2679, mul_val1_2664) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc_2606_delayed_1_0_2679, mul_val1_2664, tmp_var);
      ADD_i16_i16_2683_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2686_inst
    process(mul_val2_2670, mul_val3_2676) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val2_2670, mul_val3_2676, tmp_var);
      ADD_i16_i16_2686_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2687_inst
    process(ADD_i16_i16_2683_wire, ADD_i16_i16_2686_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i16_i16_2683_wire, ADD_i16_i16_2686_wire, tmp_var);
      acc_val_2688 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2753_inst
    process(chl_2479) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_2479, konst_2752_wire_constant, tmp_var);
      ADD_u16_u16_2753_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2773_inst
    process(col_2468) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_2468, konst_2772_wire_constant, tmp_var);
      ADD_u16_u16_2773_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2782_inst
    process(row_2463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_2463, konst_2781_wire_constant, tmp_var);
      ADD_u16_u16_2782_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u2_u2_2762_inst
    process(num_2473) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_2473, konst_2761_wire_constant, tmp_var);
      ADD_u2_u2_2762_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2552_inst
    process(ULT_u16_u1_2548_wire, UGT_u2_u1_2551_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ULT_u16_u1_2548_wire, UGT_u2_u1_2551_wire, tmp_var);
      write_input_2553 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2594_inst
    process(EQ_u16_u1_2590_wire, EQ_u16_u1_2593_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u16_u1_2590_wire, EQ_u16_u1_2593_wire, tmp_var);
      read_k_2595 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2699_inst
    process(EQ_u2_u1_2697_wire, chl_done_2693) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_2697_wire, chl_done_2693, tmp_var);
      num_done_2700 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2709_inst
    process(col_done_2705, num_done_2700) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_2705, num_done_2700, tmp_var);
      row_done_2710 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2719_inst
    process(out_done_flag_2715, col_done_2705) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2715, col_done_2705, tmp_var);
      AND_u1_u1_2719_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2725_inst
    process(out_done_flag_2715, row_done_2710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2715, row_done_2710, tmp_var);
      all_done_flag_2726 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2488_inst
    process(col_2468) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2468, konst_2487_wire_constant, tmp_var);
      EQ_u16_u1_2488_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2590_inst
    process(col_2468) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2468, konst_2589_wire_constant, tmp_var);
      EQ_u16_u1_2590_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2593_inst
    process(row_2463) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_2463, konst_2592_wire_constant, tmp_var);
      EQ_u16_u1_2593_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2692_inst
    process(chl_2479, num_chl_2454) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(chl_2479, num_chl_2454, tmp_var);
      chl_done_2693 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2704_inst
    process(col_2468, num_col_2449) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2468, num_col_2449, tmp_var);
      col_done_2705 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2714_inst
    process(row_2463, num_row_2444) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_2463, num_row_2444, tmp_var);
      out_done_flag_2715 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2491_inst
    process(num_2473) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2473, konst_2490_wire_constant, tmp_var);
      EQ_u2_u1_2491_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2697_inst
    process(num_2473) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2473, konst_2696_wire_constant, tmp_var);
      EQ_u2_u1_2697_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2662_inst
    process(kval1_2650, ival1_2578) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2650, ival1_2578, tmp_var);
      MUL_i16_i16_2662_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2668_inst
    process(kval2_2654, ival2_2582) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2654, ival2_2582, tmp_var);
      MUL_i16_i16_2668_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2674_inst
    process(kval3_2658, ival3_2586) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2658, ival3_2586, tmp_var);
      MUL_i16_i16_2674_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2720_inst
    process(AND_u1_u1_2719_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AND_u1_u1_2719_wire, tmp_var);
      store_kernel_2721 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2805_inst
    process(all_done_flag_2726) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_2726, tmp_var);
      NOT_u1_u1_2805_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2492_inst
    process(EQ_u16_u1_2488_wire, EQ_u2_u1_2491_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u16_u1_2488_wire, EQ_u2_u1_2491_wire, tmp_var);
      read_ip_2493 <= tmp_var; --
    end process;
    -- shared split operator group (27) : SUB_u16_u16_2443_inst 
    ApIntSub_group_27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2441_wire;
      num_row_2444 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2443_inst_req_0;
      SUB_u16_u16_2443_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2443_inst_req_1;
      SUB_u16_u16_2443_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_27_gI: SplitGuardInterface generic map(name => "ApIntSub_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : SUB_u16_u16_2448_inst 
    ApIntSub_group_28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2446_wire;
      num_col_2449 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2448_inst_req_0;
      SUB_u16_u16_2448_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2448_inst_req_1;
      SUB_u16_u16_2448_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_28_gI: SplitGuardInterface generic map(name => "ApIntSub_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : SUB_u16_u16_2453_inst 
    ApIntSub_group_29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_size_pipe_2451_wire;
      num_chl_2454 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2453_inst_req_0;
      SUB_u16_u16_2453_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2453_inst_req_1;
      SUB_u16_u16_2453_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_29_gI: SplitGuardInterface generic map(name => "ApIntSub_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- binary operator UGT_u2_u1_2551_inst
    process(num_2473) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_2473, konst_2550_wire_constant, tmp_var);
      UGT_u2_u1_2551_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_2548_inst
    process(col_2468, num_col_2449) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(col_2468, num_col_2449, tmp_var);
      ULT_u16_u1_2548_wire <= tmp_var; --
    end process;
    xxconvolvexxconv_ip1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip1_pipe_read_req,
        read_ack => xxconvolvexxconv_ip1_pipe_read_ack,
        read_data => xxconvolvexxconv_ip1_pipe_read_data,
        write_req => xxconvolvexxconv_ip1_pipe_write_req,
        write_ack => xxconvolvexxconv_ip1_pipe_write_ack,
        write_data => xxconvolvexxconv_ip1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip2_pipe_read_req,
        read_ack => xxconvolvexxconv_ip2_pipe_read_ack,
        read_data => xxconvolvexxconv_ip2_pipe_read_data,
        write_req => xxconvolvexxconv_ip2_pipe_write_req,
        write_ack => xxconvolvexxconv_ip2_pipe_write_ack,
        write_data => xxconvolvexxconv_ip2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip3_pipe_read_req,
        read_ack => xxconvolvexxconv_ip3_pipe_read_ack,
        read_data => xxconvolvexxconv_ip3_pipe_read_data,
        write_req => xxconvolvexxconv_ip3_pipe_write_req,
        write_ack => xxconvolvexxconv_ip3_pipe_write_ack,
        write_data => xxconvolvexxconv_ip3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k1_pipe_read_req,
        read_ack => xxconvolvexxconv_k1_pipe_read_ack,
        read_data => xxconvolvexxconv_k1_pipe_read_data,
        write_req => xxconvolvexxconv_k1_pipe_write_req,
        write_ack => xxconvolvexxconv_k1_pipe_write_ack,
        write_data => xxconvolvexxconv_k1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k2_pipe_read_req,
        read_ack => xxconvolvexxconv_k2_pipe_read_ack,
        read_data => xxconvolvexxconv_k2_pipe_read_data,
        write_req => xxconvolvexxconv_k2_pipe_write_req,
        write_ack => xxconvolvexxconv_k2_pipe_write_ack,
        write_data => xxconvolvexxconv_k2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k3_pipe_read_req,
        read_ack => xxconvolvexxconv_k3_pipe_read_ack,
        read_data => xxconvolvexxconv_k3_pipe_read_data,
        write_req => xxconvolvexxconv_k3_pipe_write_req,
        write_ack => xxconvolvexxconv_k3_pipe_write_ack,
        write_data => xxconvolvexxconv_k3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : RPIPE_input_pipe1_2496_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_2496_inst_req_0;
      RPIPE_input_pipe1_2496_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_2496_inst_req_1;
      RPIPE_input_pipe1_2496_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2493(0);
      temp2_1_2497 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_input_pipe2_2500_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe2_2500_inst_req_0;
      RPIPE_input_pipe2_2500_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe2_2500_inst_req_1;
      RPIPE_input_pipe2_2500_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2493(0);
      temp2_2_2501 <= data_out(15 downto 0);
      input_pipe2_read_1_gI: SplitGuardInterface generic map(name => "input_pipe2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe2_read_1: InputPortRevised -- 
        generic map ( name => "input_pipe2_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe2_pipe_read_req(0),
          oack => input_pipe2_pipe_read_ack(0),
          odata => input_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_input_pipe3_2504_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe3_2504_inst_req_0;
      RPIPE_input_pipe3_2504_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe3_2504_inst_req_1;
      RPIPE_input_pipe3_2504_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2493(0);
      temp2_3_2505 <= data_out(15 downto 0);
      input_pipe3_read_2_gI: SplitGuardInterface generic map(name => "input_pipe3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe3_read_2: InputPortRevised -- 
        generic map ( name => "input_pipe3_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe3_pipe_read_req(0),
          oack => input_pipe3_pipe_read_ack(0),
          odata => input_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_kernel_pipe1_2598_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_2598_inst_req_0;
      RPIPE_kernel_pipe1_2598_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_2598_inst_req_1;
      RPIPE_kernel_pipe1_2598_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2595(0);
      tempk1_1_2599 <= data_out(15 downto 0);
      kernel_pipe1_read_3_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_3: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_kernel_pipe2_2602_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_2602_inst_req_0;
      RPIPE_kernel_pipe2_2602_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_2602_inst_req_1;
      RPIPE_kernel_pipe2_2602_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2595(0);
      tempk1_2_2603 <= data_out(15 downto 0);
      kernel_pipe2_read_4_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_4: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_4", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : RPIPE_kernel_pipe3_2606_inst 
    InportGroup_5: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe3_2606_inst_req_0;
      RPIPE_kernel_pipe3_2606_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe3_2606_inst_req_1;
      RPIPE_kernel_pipe3_2606_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2595(0);
      tempk1_3_2607 <= data_out(15 downto 0);
      kernel_pipe3_read_5_gI: SplitGuardInterface generic map(name => "kernel_pipe3_read_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_read_5: InputPortRevised -- 
        generic map ( name => "kernel_pipe3_read_5", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe3_pipe_read_req(0),
          oack => kernel_pipe3_pipe_read_ack(0),
          odata => kernel_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : RPIPE_num_out_pipe_2441_inst RPIPE_num_out_pipe_2446_inst 
    InportGroup_6: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_num_out_pipe_2441_inst_req_0;
      reqL_unguarded(0) <= RPIPE_num_out_pipe_2446_inst_req_0;
      RPIPE_num_out_pipe_2441_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_num_out_pipe_2446_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_num_out_pipe_2441_inst_req_1;
      reqR_unguarded(0) <= RPIPE_num_out_pipe_2446_inst_req_1;
      RPIPE_num_out_pipe_2441_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_num_out_pipe_2446_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      RPIPE_num_out_pipe_2441_wire <= data_out(31 downto 16);
      RPIPE_num_out_pipe_2446_wire <= data_out(15 downto 0);
      num_out_pipe_read_6_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_6_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_6: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_6", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : RPIPE_size_pipe_2451_inst 
    InportGroup_7: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_2451_inst_req_0;
      RPIPE_size_pipe_2451_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_2451_inst_req_1;
      RPIPE_size_pipe_2451_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_size_pipe_2451_wire <= data_out(15 downto 0);
      size_pipe_read_7_gI: SplitGuardInterface generic map(name => "size_pipe_read_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_7: InputPortRevised -- 
        generic map ( name => "size_pipe_read_7", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : RPIPE_xxconvolvexxconv_ip1_2508_inst 
    InportGroup_8: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2508_inst_req_0;
      RPIPE_xxconvolvexxconv_ip1_2508_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2508_inst_req_1;
      RPIPE_xxconvolvexxconv_ip1_2508_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2493(0);
      temp1_1_2509 <= data_out(15 downto 0);
      xxconvolvexxconv_ip1_read_8_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_read_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_read_8: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1_read_8", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip1_pipe_read_req(0),
          oack => xxconvolvexxconv_ip1_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : RPIPE_xxconvolvexxconv_ip2_2512_inst 
    InportGroup_9: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2512_inst_req_0;
      RPIPE_xxconvolvexxconv_ip2_2512_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2512_inst_req_1;
      RPIPE_xxconvolvexxconv_ip2_2512_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2493(0);
      temp1_2_2513 <= data_out(15 downto 0);
      xxconvolvexxconv_ip2_read_9_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_read_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_read_9: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2_read_9", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip2_pipe_read_req(0),
          oack => xxconvolvexxconv_ip2_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : RPIPE_xxconvolvexxconv_ip3_2516_inst 
    InportGroup_10: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2516_inst_req_0;
      RPIPE_xxconvolvexxconv_ip3_2516_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2516_inst_req_1;
      RPIPE_xxconvolvexxconv_ip3_2516_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2493(0);
      temp1_3_2517 <= data_out(15 downto 0);
      xxconvolvexxconv_ip3_read_10_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_read_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_read_10: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3_read_10", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip3_pipe_read_req(0),
          oack => xxconvolvexxconv_ip3_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : RPIPE_xxconvolvexxconv_k1_2610_inst 
    InportGroup_11: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2610_inst_req_0;
      RPIPE_xxconvolvexxconv_k1_2610_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2610_inst_req_1;
      RPIPE_xxconvolvexxconv_k1_2610_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2595(0);
      tempk2_1_2611 <= data_out(15 downto 0);
      xxconvolvexxconv_k1_read_11_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_read_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_read_11: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1_read_11", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k1_pipe_read_req(0),
          oack => xxconvolvexxconv_k1_pipe_read_ack(0),
          odata => xxconvolvexxconv_k1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- shared inport operator group (12) : RPIPE_xxconvolvexxconv_k2_2614_inst 
    InportGroup_12: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2614_inst_req_0;
      RPIPE_xxconvolvexxconv_k2_2614_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2614_inst_req_1;
      RPIPE_xxconvolvexxconv_k2_2614_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2595(0);
      tempk2_2_2615 <= data_out(15 downto 0);
      xxconvolvexxconv_k2_read_12_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_read_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_read_12: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2_read_12", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k2_pipe_read_req(0),
          oack => xxconvolvexxconv_k2_pipe_read_ack(0),
          odata => xxconvolvexxconv_k2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 12
    -- shared inport operator group (13) : RPIPE_xxconvolvexxconv_k3_2618_inst 
    InportGroup_13: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2618_inst_req_0;
      RPIPE_xxconvolvexxconv_k3_2618_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2618_inst_req_1;
      RPIPE_xxconvolvexxconv_k3_2618_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2595(0);
      tempk2_3_2619 <= data_out(15 downto 0);
      xxconvolvexxconv_k3_read_13_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_read_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_read_13: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3_read_13", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k3_pipe_read_req(0),
          oack => xxconvolvexxconv_k3_pipe_read_ack(0),
          odata => xxconvolvexxconv_k3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 13
    -- shared outport operator group (0) : WPIPE_input_done_pipe_2806_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_2806_inst_req_0;
      WPIPE_input_done_pipe_2806_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_2806_inst_req_1;
      WPIPE_input_done_pipe_2806_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2807_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_output_pipe_2799_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_output_pipe_2799_inst_req_0;
      WPIPE_output_pipe_2799_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_output_pipe_2799_inst_req_1;
      WPIPE_output_pipe_2799_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= num_done_2708_delayed_1_0_2797(0);
      data_in <= type_cast_2801_wire;
      output_pipe_write_1_gI: SplitGuardInterface generic map(name => "output_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_xxconvolvexxconv_ip1_2558_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2558_inst_req_0;
      WPIPE_xxconvolvexxconv_ip1_2558_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2558_inst_req_1;
      WPIPE_xxconvolvexxconv_ip1_2558_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2500_delayed_1_0_2556(0);
      data_in <= iread1_2526;
      xxconvolvexxconv_ip1_write_2_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_write_2: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip1_pipe_write_req(0),
          oack => xxconvolvexxconv_ip1_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_xxconvolvexxconv_ip2_2565_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2565_inst_req_0;
      WPIPE_xxconvolvexxconv_ip2_2565_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2565_inst_req_1;
      WPIPE_xxconvolvexxconv_ip2_2565_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2504_delayed_1_0_2563(0);
      data_in <= iread2_2535;
      xxconvolvexxconv_ip2_write_3_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_write_3: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip2_pipe_write_req(0),
          oack => xxconvolvexxconv_ip2_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_xxconvolvexxconv_ip3_2572_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2572_inst_req_0;
      WPIPE_xxconvolvexxconv_ip3_2572_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2572_inst_req_1;
      WPIPE_xxconvolvexxconv_ip3_2572_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2508_delayed_1_0_2570(0);
      data_in <= iread3_2544;
      xxconvolvexxconv_ip3_write_4_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_write_4: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip3_pipe_write_req(0),
          oack => xxconvolvexxconv_ip3_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_xxconvolvexxconv_k1_2731_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2731_inst_req_0;
      WPIPE_xxconvolvexxconv_k1_2731_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2731_inst_req_1;
      WPIPE_xxconvolvexxconv_k1_2731_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2652_delayed_1_0_2729(0);
      data_in <= kread1_2628;
      xxconvolvexxconv_k1_write_5_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_write_5: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k1_pipe_write_req(0),
          oack => xxconvolvexxconv_k1_pipe_write_ack(0),
          odata => xxconvolvexxconv_k1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_xxconvolvexxconv_k2_2738_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2738_inst_req_0;
      WPIPE_xxconvolvexxconv_k2_2738_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2738_inst_req_1;
      WPIPE_xxconvolvexxconv_k2_2738_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2656_delayed_1_0_2736(0);
      data_in <= kread2_2637;
      xxconvolvexxconv_k2_write_6_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_write_6: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k2_pipe_write_req(0),
          oack => xxconvolvexxconv_k2_pipe_write_ack(0),
          odata => xxconvolvexxconv_k2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_xxconvolvexxconv_k3_2745_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2745_inst_req_0;
      WPIPE_xxconvolvexxconv_k3_2745_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2745_inst_req_1;
      WPIPE_xxconvolvexxconv_k3_2745_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2660_delayed_1_0_2743(0);
      data_in <= kread3_2646;
      xxconvolvexxconv_k3_write_7_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_write_7: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k3_pipe_write_req(0),
          oack => xxconvolvexxconv_k3_pipe_write_ack(0),
          odata => xxconvolvexxconv_k3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    num_chl : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal num_chl_buffer :  std_logic_vector(15 downto 0);
  signal num_chl_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_1309_start: Boolean;
  signal loadKernelChannel_CP_1309_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_410_index_offset_ack_0 : boolean;
  signal nfetch_val_543_455_buf_ack_0 : boolean;
  signal ptr_deref_415_load_0_ack_0 : boolean;
  signal addr_of_411_final_reg_ack_1 : boolean;
  signal ptr_deref_415_load_0_ack_1 : boolean;
  signal array_obj_ref_410_index_offset_ack_1 : boolean;
  signal array_obj_ref_410_index_offset_req_1 : boolean;
  signal nmycount_471_452_buf_ack_1 : boolean;
  signal start_add_451_buf_ack_0 : boolean;
  signal phi_stmt_453_ack_0 : boolean;
  signal my_fetch_416_456_buf_req_0 : boolean;
  signal array_obj_ref_410_index_offset_req_0 : boolean;
  signal RPIPE_input_done_pipe_444_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_444_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_444_inst_ack_0 : boolean;
  signal nfetch_val_543_455_buf_ack_1 : boolean;
  signal RPIPE_input_done_pipe_444_inst_req_0 : boolean;
  signal nfetch_val_543_455_buf_req_0 : boolean;
  signal phi_stmt_449_ack_0 : boolean;
  signal nfetch_val_543_455_buf_req_1 : boolean;
  signal phi_stmt_449_req_0 : boolean;
  signal start_add_451_buf_ack_1 : boolean;
  signal ptr_deref_415_load_0_req_1 : boolean;
  signal start_add_451_buf_req_1 : boolean;
  signal phi_stmt_453_req_1 : boolean;
  signal addr_of_411_final_reg_req_1 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_ack_1 : boolean;
  signal do_while_stmt_447_branch_req_0 : boolean;
  signal start_add_451_buf_req_0 : boolean;
  signal my_fetch_416_456_buf_ack_1 : boolean;
  signal WPIPE_kernel_pipe3_505_inst_req_1 : boolean;
  signal nmycount_471_452_buf_req_0 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_req_0 : boolean;
  signal nmycount_471_452_buf_ack_0 : boolean;
  signal my_fetch_416_456_buf_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_501_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_505_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe3_505_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_501_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_505_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe2_501_inst_ack_1 : boolean;
  signal addr_of_411_final_reg_ack_0 : boolean;
  signal phi_stmt_453_req_0 : boolean;
  signal ptr_deref_415_load_0_req_0 : boolean;
  signal phi_stmt_449_req_1 : boolean;
  signal my_fetch_416_456_buf_req_1 : boolean;
  signal nmycount_471_452_buf_req_1 : boolean;
  signal WPIPE_kernel_pipe2_501_inst_ack_0 : boolean;
  signal addr_of_411_final_reg_req_0 : boolean;
  signal array_obj_ref_521_index_offset_req_0 : boolean;
  signal array_obj_ref_521_index_offset_ack_0 : boolean;
  signal array_obj_ref_521_index_offset_req_1 : boolean;
  signal array_obj_ref_521_index_offset_ack_1 : boolean;
  signal addr_of_522_final_reg_req_0 : boolean;
  signal addr_of_522_final_reg_ack_0 : boolean;
  signal addr_of_522_final_reg_req_1 : boolean;
  signal addr_of_522_final_reg_ack_1 : boolean;
  signal W_fn_488_delayed_7_0_524_inst_req_0 : boolean;
  signal W_fn_488_delayed_7_0_524_inst_ack_0 : boolean;
  signal W_fn_488_delayed_7_0_524_inst_req_1 : boolean;
  signal W_fn_488_delayed_7_0_524_inst_ack_1 : boolean;
  signal ptr_deref_530_load_0_req_0 : boolean;
  signal ptr_deref_530_load_0_ack_0 : boolean;
  signal ptr_deref_530_load_0_req_1 : boolean;
  signal ptr_deref_530_load_0_ack_1 : boolean;
  signal W_fn_494_delayed_13_0_532_inst_req_0 : boolean;
  signal W_fn_494_delayed_13_0_532_inst_ack_0 : boolean;
  signal W_fn_494_delayed_13_0_532_inst_req_1 : boolean;
  signal W_fn_494_delayed_13_0_532_inst_ack_1 : boolean;
  signal W_fetch_val_496_delayed_13_0_535_inst_req_0 : boolean;
  signal W_fetch_val_496_delayed_13_0_535_inst_ack_0 : boolean;
  signal W_fetch_val_496_delayed_13_0_535_inst_req_1 : boolean;
  signal W_fetch_val_496_delayed_13_0_535_inst_ack_1 : boolean;
  signal do_while_stmt_447_branch_ack_0 : boolean;
  signal do_while_stmt_447_branch_ack_1 : boolean;
  signal WPIPE_size_pipe_551_inst_req_0 : boolean;
  signal WPIPE_size_pipe_551_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_551_inst_req_1 : boolean;
  signal WPIPE_size_pipe_551_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(79 downto 64) <= num_chl;
  num_chl_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_1309_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1309_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1309_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1309_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_1309: Block -- control-path 
    signal loadKernelChannel_CP_1309_elements: BooleanArray(98 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_1309_elements(0) <= loadKernelChannel_CP_1309_start;
    loadKernelChannel_CP_1309_symbol <= loadKernelChannel_CP_1309_elements(98);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Sample/rr
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_computed_1
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_index_resized_1
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_sample_start_
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_update_start_
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_complete/req
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/$entry
      -- CP-element group 0: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_complete/$entry
      -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => addr_of_411_final_reg_req_1); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => array_obj_ref_410_index_offset_req_0); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => array_obj_ref_410_index_offset_req_1); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => ptr_deref_415_load_0_req_1); -- 
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => RPIPE_input_done_pipe_444_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Sample/ack
      -- CP-element group 1: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_sample_complete
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_index_offset_ack_0, ack => loadKernelChannel_CP_1309_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_sample_start_
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_request/$entry
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_offset_calculated
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/array_obj_ref_410_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_request/req
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_index_offset_ack_1, ack => loadKernelChannel_CP_1309_elements(2)); -- 
    req_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(2), ack => addr_of_411_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_sample_completed_
      -- CP-element group 3: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_request/ack
      -- CP-element group 3: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_request/$exit
      -- 
    ack_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_411_final_reg_ack_0, ack => loadKernelChannel_CP_1309_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_sample_start_
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_complete/ack
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_address_resized
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_update_completed_
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/addr_of_411_complete/$exit
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/word_access_start/word_0/rr
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_411_final_reg_ack_1, ack => loadKernelChannel_CP_1309_elements(4)); -- 
    rr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(4), ack => ptr_deref_415_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_sample_completed_
      -- CP-element group 5: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Sample/$exit
      -- 
    ra_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_415_load_0_ack_0, ack => loadKernelChannel_CP_1309_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/ptr_deref_415_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/ptr_deref_415_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_update_completed_
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/ptr_deref_415_Merge/merge_ack
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/ptr_deref_415_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_400_to_assign_stmt_445/ptr_deref_415_Update/$exit
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_415_load_0_ack_1, ack => loadKernelChannel_CP_1309_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Update/cr
      -- CP-element group 7: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Update/$entry
      -- CP-element group 7: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Sample/ra
      -- CP-element group 7: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_update_start_
      -- CP-element group 7: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_sample_completed_
      -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_444_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(7)); -- 
    cr_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(7), ack => RPIPE_input_done_pipe_444_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Update/ca
      -- CP-element group 8: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_Update/$exit
      -- CP-element group 8: 	 assign_stmt_400_to_assign_stmt_445/RPIPE_input_done_pipe_444_update_completed_
      -- 
    ca_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_444_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_446/do_while_stmt_447__entry__
      -- CP-element group 9: 	 branch_block_stmt_446/$entry
      -- CP-element group 9: 	 assign_stmt_400_to_assign_stmt_445/$exit
      -- CP-element group 9: 	 branch_block_stmt_446/branch_block_stmt_446__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(1) & loadKernelChannel_CP_1309_elements(6) & loadKernelChannel_CP_1309_elements(8);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	96 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	97 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_446/do_while_stmt_447__exit__
      -- CP-element group 10: 	 branch_block_stmt_446/$exit
      -- CP-element group 10: 	 branch_block_stmt_446/branch_block_stmt_446__exit__
      -- CP-element group 10: 	 assign_stmt_553/$entry
      -- CP-element group 10: 	 assign_stmt_553/WPIPE_size_pipe_551_sample_start_
      -- CP-element group 10: 	 assign_stmt_553/WPIPE_size_pipe_551_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_553/WPIPE_size_pipe_551_Sample/req
      -- 
    req_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(10), ack => WPIPE_size_pipe_551_inst_req_0); -- 
    loadKernelChannel_CP_1309_elements(10) <= loadKernelChannel_CP_1309_elements(96);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_446/do_while_stmt_447/$entry
      -- CP-element group 11: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447__entry__
      -- 
    loadKernelChannel_CP_1309_elements(11) <= loadKernelChannel_CP_1309_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	96 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447__exit__
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_446/do_while_stmt_447/loop_back
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	94 
    -- CP-element group 14: 	95 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_446/do_while_stmt_447/condition_done
      -- CP-element group 14: 	 branch_block_stmt_446/do_while_stmt_447/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_446/do_while_stmt_447/loop_taken/$entry
      -- 
    loadKernelChannel_CP_1309_elements(14) <= loadKernelChannel_CP_1309_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	93 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_446/do_while_stmt_447/loop_body_done
      -- 
    loadKernelChannel_CP_1309_elements(15) <= loadKernelChannel_CP_1309_elements(93);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_1309_elements(16) <= loadKernelChannel_CP_1309_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_1309_elements(17) <= loadKernelChannel_CP_1309_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	70 
    -- CP-element group 18: 	71 
    -- CP-element group 18: 	92 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	27 
    -- CP-element group 19: 	92 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/condition_evaluated
      -- 
    condition_evaluated_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(19), ack => do_while_stmt_447_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(23) & loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(92);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	41 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/aggregated_phi_sample_req
      -- CP-element group 20: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_sample_start__ps
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(24) & loadKernelChannel_CP_1309_elements(41) & loadKernelChannel_CP_1309_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	81 
    -- CP-element group 21: 	85 
    -- CP-element group 21: 	89 
    -- CP-element group 21: 	93 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	41 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/aggregated_phi_sample_ack
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(26) & loadKernelChannel_CP_1309_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/aggregated_phi_update_req
      -- CP-element group 22: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_update_start__ps
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(25) & loadKernelChannel_CP_1309_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	64 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	78 
    -- CP-element group 25: 	86 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(61) & loadKernelChannel_CP_1309_elements(64) & loadKernelChannel_CP_1309_elements(67) & loadKernelChannel_CP_1309_elements(72) & loadKernelChannel_CP_1309_elements(78) & loadKernelChannel_CP_1309_elements(86);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	60 
    -- CP-element group 27: 	63 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	72 
    -- CP-element group 27: 	76 
    -- CP-element group 27: 	84 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Sample/req
      -- 
    req_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(27), ack => array_obj_ref_521_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_loopback_trigger
      -- 
    loadKernelChannel_CP_1309_elements(28) <= loadKernelChannel_CP_1309_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_loopback_sample_req_ps
      -- CP-element group 29: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_loopback_sample_req
      -- 
    phi_stmt_449_loopback_sample_req_1461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_449_loopback_sample_req_1461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(29), ack => phi_stmt_449_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_entry_trigger
      -- 
    loadKernelChannel_CP_1309_elements(30) <= loadKernelChannel_CP_1309_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_entry_sample_req_ps
      -- CP-element group 31: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_entry_sample_req
      -- 
    phi_stmt_449_entry_sample_req_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_449_entry_sample_req_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(31), ack => phi_stmt_449_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_phi_mux_ack_ps
      -- CP-element group 32: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_449_phi_mux_ack
      -- 
    phi_stmt_449_phi_mux_ack_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_449_ack_0, ack => loadKernelChannel_CP_1309_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Sample/req
      -- CP-element group 33: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Sample/$entry
      -- 
    req_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(33), ack => start_add_451_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_update_start_
      -- CP-element group 34: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Update/req
      -- 
    req_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(34), ack => start_add_451_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Sample/$exit
      -- 
    ack_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_451_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_start_add_451_update_completed_
      -- 
    ack_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_451_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_sample_start__ps
      -- CP-element group 37: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Sample/req
      -- 
    req_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(37), ack => nmycount_471_452_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_update_start_
      -- CP-element group 38: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Update/req
      -- 
    req_1503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(38), ack => nmycount_471_452_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Sample/ack
      -- 
    ack_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_471_452_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nmycount_452_Update/$exit
      -- 
    ack_1504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_471_452_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	21 
    -- CP-element group 41: 	83 
    -- CP-element group 41: 	87 
    -- CP-element group 41: 	91 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(83) & loadKernelChannel_CP_1309_elements(87) & loadKernelChannel_CP_1309_elements(91);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	64 
    -- CP-element group 42: 	67 
    -- CP-element group 42: 	90 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(61) & loadKernelChannel_CP_1309_elements(64) & loadKernelChannel_CP_1309_elements(67) & loadKernelChannel_CP_1309_elements(90);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_sample_start__ps
      -- 
    loadKernelChannel_CP_1309_elements(43) <= loadKernelChannel_CP_1309_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_update_start__ps
      -- 
    loadKernelChannel_CP_1309_elements(45) <= loadKernelChannel_CP_1309_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	63 
    -- CP-element group 46: 	66 
    -- CP-element group 46: 	88 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_update_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_loopback_trigger
      -- 
    loadKernelChannel_CP_1309_elements(47) <= loadKernelChannel_CP_1309_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_loopback_sample_req
      -- CP-element group 48: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_loopback_sample_req_ps
      -- 
    phi_stmt_453_loopback_sample_req_1515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_loopback_sample_req_1515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(48), ack => phi_stmt_453_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_entry_trigger
      -- 
    loadKernelChannel_CP_1309_elements(49) <= loadKernelChannel_CP_1309_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_entry_sample_req_ps
      -- CP-element group 50: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_entry_sample_req
      -- 
    phi_stmt_453_entry_sample_req_1518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_entry_sample_req_1518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(50), ack => phi_stmt_453_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_phi_mux_ack_ps
      -- CP-element group 51: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/phi_stmt_453_phi_mux_ack
      -- 
    phi_stmt_453_phi_mux_ack_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_453_ack_0, ack => loadKernelChannel_CP_1309_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Sample/req
      -- 
    req_1534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(52), ack => nfetch_val_543_455_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Update/req
      -- CP-element group 53: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_update_start_
      -- 
    req_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(53), ack => nfetch_val_543_455_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Sample/$exit
      -- 
    ack_1535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_543_455_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_nfetch_val_455_update_completed_
      -- 
    ack_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_543_455_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_sample_start_
      -- 
    req_1552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(56), ack => my_fetch_416_456_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_update_start_
      -- CP-element group 57: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Update/req
      -- 
    req_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(57), ack => my_fetch_416_456_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_sample_completed__ps
      -- 
    ack_1553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_416_456_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/R_my_fetch_456_update_completed__ps
      -- 
    ack_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_416_456_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_sample_start_
      -- 
    req_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(60), ack => WPIPE_kernel_pipe1_497_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Update/req
      -- CP-element group 61: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_update_start_
      -- CP-element group 61: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_sample_completed_
      -- 
    ack_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_497_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(61)); -- 
    req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(61), ack => WPIPE_kernel_pipe1_497_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	93 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe1_497_update_completed_
      -- 
    ack_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_497_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	27 
    -- CP-element group 63: 	46 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Sample/req
      -- 
    req_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(63), ack => WPIPE_kernel_pipe2_501_inst_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(65);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	25 
    -- CP-element group 64: 	42 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_update_start_
      -- CP-element group 64: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Update/req
      -- CP-element group 64: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Sample/ack
      -- 
    ack_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_501_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(64)); -- 
    req_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(64), ack => WPIPE_kernel_pipe2_501_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	93 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe2_501_Update/ack
      -- 
    ack_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_501_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: 	46 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Sample/req
      -- CP-element group 66: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Sample/$entry
      -- 
    req_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(66), ack => WPIPE_kernel_pipe3_505_inst_req_0); -- 
    loadKernelChannel_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(68);
      gj_loadKernelChannel_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	42 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Update/req
      -- CP-element group 67: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_update_start_
      -- CP-element group 67: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Sample/$exit
      -- 
    ack_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_505_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(67)); -- 
    req_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(67), ack => WPIPE_kernel_pipe3_505_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	93 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/WPIPE_kernel_pipe3_505_Update/ack
      -- 
    ack_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_505_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	73 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_request/$entry
      -- CP-element group 69: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_request/req
      -- 
    req_1641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(69), ack => addr_of_522_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(73) & loadKernelChannel_CP_1309_elements(74);
      gj_loadKernelChannel_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	18 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	75 
    -- CP-element group 70: 	82 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	75 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_update_start_
      -- CP-element group 70: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_complete/$entry
      -- CP-element group 70: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_complete/req
      -- 
    req_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(70), ack => addr_of_522_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(75) & loadKernelChannel_CP_1309_elements(82);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	18 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	74 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_update_start
      -- CP-element group 71: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Update/req
      -- 
    req_1631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(71), ack => array_obj_ref_521_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(73) & loadKernelChannel_CP_1309_elements(74);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	27 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	93 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_sample_complete
      -- CP-element group 72: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Sample/ack
      -- 
    ack_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_521_index_offset_ack_0, ack => loadKernelChannel_CP_1309_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (8) 
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_offset_calculated
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_final_index_sum_regn_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/array_obj_ref_521_base_plus_offset/sum_rename_ack
      -- 
    ack_1632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_521_index_offset_ack_1, ack => loadKernelChannel_CP_1309_elements(73)); -- 
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	71 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_request/$exit
      -- CP-element group 74: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_request/ack
      -- 
    ack_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_522_final_reg_ack_0, ack => loadKernelChannel_CP_1309_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	70 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	80 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	70 
    -- CP-element group 75:  members (19) 
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_word_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/addr_of_522_complete/ack
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_root_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_address_resized
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_addr_resize/$entry
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_addr_resize/$exit
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_addr_resize/base_resize_req
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_addr_resize/base_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_plus_offset/$entry
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_plus_offset/$exit
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_plus_offset/sum_rename_req
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_base_plus_offset/sum_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_word_addrgen/$entry
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_word_addrgen/$exit
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_word_addrgen/root_register_req
      -- CP-element group 75: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_word_addrgen/root_register_ack
      -- 
    ack_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_522_final_reg_ack_1, ack => loadKernelChannel_CP_1309_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	27 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Sample/req
      -- 
    req_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(76), ack => W_fn_488_delayed_7_0_524_inst_req_0); -- 
    loadKernelChannel_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(78);
      gj_loadKernelChannel_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	82 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_update_start_
      -- CP-element group 77: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Update/req
      -- 
    req_1660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(77), ack => W_fn_488_delayed_7_0_524_inst_req_1); -- 
    loadKernelChannel_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(79) & loadKernelChannel_CP_1309_elements(82);
      gj_loadKernelChannel_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	25 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Sample/ack
      -- 
    ack_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_488_delayed_7_0_524_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_526_Update/ack
      -- 
    ack_1661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_488_delayed_7_0_524_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: 	79 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/word_access_start/word_0/rr
      -- 
    rr_1694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(80), ack => ptr_deref_530_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(75) & loadKernelChannel_CP_1309_elements(79) & loadKernelChannel_CP_1309_elements(82);
      gj_loadKernelChannel_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	21 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_update_start_
      -- CP-element group 81: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/word_access_complete/word_0/cr
      -- 
    cr_1705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(81), ack => ptr_deref_530_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(83);
      gj_loadKernelChannel_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/word_access_start/$exit
      -- CP-element group 82: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Sample/word_access_start/word_0/ra
      -- 
    ra_1695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_530_load_0_ack_0, ack => loadKernelChannel_CP_1309_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	93 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	41 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/word_access_complete/$exit
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/word_access_complete/word_0/ca
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/ptr_deref_530_Merge/$entry
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/ptr_deref_530_Merge/$exit
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/ptr_deref_530_Merge/merge_req
      -- CP-element group 83: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/ptr_deref_530_Update/ptr_deref_530_Merge/merge_ack
      -- 
    ca_1706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_530_load_0_ack_1, ack => loadKernelChannel_CP_1309_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	27 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Sample/req
      -- 
    req_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(84), ack => W_fn_494_delayed_13_0_532_inst_req_0); -- 
    loadKernelChannel_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(86);
      gj_loadKernelChannel_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	21 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_update_start_
      -- CP-element group 85: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Update/req
      -- 
    req_1724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(85), ack => W_fn_494_delayed_13_0_532_inst_req_1); -- 
    loadKernelChannel_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(87);
      gj_loadKernelChannel_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Sample/ack
      -- 
    ack_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_494_delayed_13_0_532_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	93 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_534_Update/ack
      -- 
    ack_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_494_delayed_13_0_532_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	46 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Sample/req
      -- 
    req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(88), ack => W_fetch_val_496_delayed_13_0_535_inst_req_0); -- 
    loadKernelChannel_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(90);
      gj_loadKernelChannel_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	21 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_update_start_
      -- CP-element group 89: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Update/req
      -- 
    req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(89), ack => W_fetch_val_496_delayed_13_0_535_inst_req_1); -- 
    loadKernelChannel_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(91);
      gj_loadKernelChannel_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	42 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Sample/ack
      -- 
    ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_496_delayed_13_0_535_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	41 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/assign_stmt_537_Update/ack
      -- 
    ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_496_delayed_13_0_535_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(91)); -- 
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	18 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	19 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_1309_elements(18), ack => loadKernelChannel_CP_1309_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	21 
    -- CP-element group 93: 	62 
    -- CP-element group 93: 	65 
    -- CP-element group 93: 	68 
    -- CP-element group 93: 	72 
    -- CP-element group 93: 	83 
    -- CP-element group 93: 	87 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	15 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_446/do_while_stmt_447/do_while_stmt_447_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(62) & loadKernelChannel_CP_1309_elements(65) & loadKernelChannel_CP_1309_elements(68) & loadKernelChannel_CP_1309_elements(72) & loadKernelChannel_CP_1309_elements(83) & loadKernelChannel_CP_1309_elements(87) & loadKernelChannel_CP_1309_elements(91);
      gj_loadKernelChannel_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_446/do_while_stmt_447/loop_exit/$exit
      -- CP-element group 94: 	 branch_block_stmt_446/do_while_stmt_447/loop_exit/ack
      -- 
    ack_1744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_447_branch_ack_0, ack => loadKernelChannel_CP_1309_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	14 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_446/do_while_stmt_447/loop_taken/$exit
      -- CP-element group 95: 	 branch_block_stmt_446/do_while_stmt_447/loop_taken/ack
      -- 
    ack_1748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_447_branch_ack_1, ack => loadKernelChannel_CP_1309_elements(95)); -- 
    -- CP-element group 96:  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	12 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	10 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_446/do_while_stmt_447/$exit
      -- 
    loadKernelChannel_CP_1309_elements(96) <= loadKernelChannel_CP_1309_elements(12);
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	10 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 assign_stmt_553/WPIPE_size_pipe_551_sample_completed_
      -- CP-element group 97: 	 assign_stmt_553/WPIPE_size_pipe_551_update_start_
      -- CP-element group 97: 	 assign_stmt_553/WPIPE_size_pipe_551_Sample/$exit
      -- CP-element group 97: 	 assign_stmt_553/WPIPE_size_pipe_551_Sample/ack
      -- CP-element group 97: 	 assign_stmt_553/WPIPE_size_pipe_551_Update/$entry
      -- CP-element group 97: 	 assign_stmt_553/WPIPE_size_pipe_551_Update/req
      -- 
    ack_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_551_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(97)); -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(97), ack => WPIPE_size_pipe_551_inst_req_1); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 $exit
      -- CP-element group 98: 	 assign_stmt_553/$exit
      -- CP-element group 98: 	 assign_stmt_553/WPIPE_size_pipe_551_update_completed_
      -- CP-element group 98: 	 assign_stmt_553/WPIPE_size_pipe_551_Update/$exit
      -- CP-element group 98: 	 assign_stmt_553/WPIPE_size_pipe_551_Update/ack
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_551_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(98)); -- 
    loadKernelChannel_do_while_stmt_447_terminator_1749: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_447_terminator_1749", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_1309_elements(15),loop_continue => loadKernelChannel_CP_1309_elements(95),loop_terminate => loadKernelChannel_CP_1309_elements(94),loop_back => loadKernelChannel_CP_1309_elements(13),loop_exit => loadKernelChannel_CP_1309_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_449_phi_seq_1505_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1309_elements(30);
      loadKernelChannel_CP_1309_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1309_elements(35);
      loadKernelChannel_CP_1309_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1309_elements(36);
      loadKernelChannel_CP_1309_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1309_elements(28);
      loadKernelChannel_CP_1309_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1309_elements(39);
      loadKernelChannel_CP_1309_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1309_elements(40);
      loadKernelChannel_CP_1309_elements(29) <= phi_mux_reqs(1);
      phi_stmt_449_phi_seq_1505 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_449_phi_seq_1505") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1309_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_1309_elements(26), 
          phi_update_req => loadKernelChannel_CP_1309_elements(22), 
          phi_update_ack => loadKernelChannel_CP_1309_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_1309_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_453_phi_seq_1559_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1309_elements(47);
      loadKernelChannel_CP_1309_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1309_elements(54);
      loadKernelChannel_CP_1309_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1309_elements(55);
      loadKernelChannel_CP_1309_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1309_elements(49);
      loadKernelChannel_CP_1309_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1309_elements(58);
      loadKernelChannel_CP_1309_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1309_elements(59);
      loadKernelChannel_CP_1309_elements(50) <= phi_mux_reqs(1);
      phi_stmt_453_phi_seq_1559 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_453_phi_seq_1559") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1309_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_1309_elements(44), 
          phi_update_req => loadKernelChannel_CP_1309_elements(45), 
          phi_update_ack => loadKernelChannel_CP_1309_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_1309_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1447_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_1309_elements(16);
        preds(1)  <= loadKernelChannel_CP_1309_elements(17);
        entry_tmerge_1447 : transition_merge -- 
          generic map(name => " entry_tmerge_1447")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_462_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_511_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_475_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_520_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_520_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_520_wire : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_485_wire : std_logic_vector(0 downto 0);
    signal R_sh_start_409_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_409_scaled : std_logic_vector(13 downto 0);
    signal SHL_u16_u16_398_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_427_wire : std_logic_vector(15 downto 0);
    signal SUB_u64_u64_463_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_548_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_488_wire : std_logic_vector(0 downto 0);
    signal ULT_u64_u1_549_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_410_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_410_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_410_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_410_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_410_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_410_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_521_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_521_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_521_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_521_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_521_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_521_root_address : std_logic_vector(13 downto 0);
    signal ea1_422 : std_logic_vector(63 downto 0);
    signal ea2_430 : std_logic_vector(63 downto 0);
    signal ea3_436 : std_logic_vector(63 downto 0);
    signal fetch_addr_412 : std_logic_vector(31 downto 0);
    signal fetch_addr_523 : std_logic_vector(31 downto 0);
    signal fetch_val_453 : std_logic_vector(63 downto 0);
    signal fetch_val_496_delayed_13_0_537 : std_logic_vector(63 downto 0);
    signal first_fill_441 : std_logic_vector(0 downto 0);
    signal fn_488_delayed_7_0_526 : std_logic_vector(0 downto 0);
    signal fn_494_delayed_13_0_534 : std_logic_vector(0 downto 0);
    signal fn_514 : std_logic_vector(0 downto 0);
    signal fv_531 : std_logic_vector(63 downto 0);
    signal konst_397_wire_constant : std_logic_vector(15 downto 0);
    signal konst_403_wire_constant : std_logic_vector(63 downto 0);
    signal konst_426_wire_constant : std_logic_vector(15 downto 0);
    signal konst_439_wire_constant : std_logic_vector(63 downto 0);
    signal konst_459_wire_constant : std_logic_vector(63 downto 0);
    signal konst_461_wire_constant : std_logic_vector(63 downto 0);
    signal konst_464_wire_constant : std_logic_vector(63 downto 0);
    signal konst_469_wire_constant : std_logic_vector(63 downto 0);
    signal konst_510_wire_constant : std_logic_vector(63 downto 0);
    signal konst_512_wire_constant : std_logic_vector(63 downto 0);
    signal konst_519_wire_constant : std_logic_vector(63 downto 0);
    signal konst_547_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_416 : std_logic_vector(63 downto 0);
    signal my_fetch_416_456_buffered : std_logic_vector(63 downto 0);
    signal my_num1_466 : std_logic_vector(63 downto 0);
    signal mycount_449 : std_logic_vector(63 downto 0);
    signal nfetch_val_543 : std_logic_vector(63 downto 0);
    signal nfetch_val_543_455_buffered : std_logic_vector(63 downto 0);
    signal nmycount_471 : std_logic_vector(63 downto 0);
    signal nmycount_471_452_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_415_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_415_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_415_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_415_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_415_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_530_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_530_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_530_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_530_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_530_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_size_400 : std_logic_vector(15 downto 0);
    signal send_to_1_482 : std_logic_vector(0 downto 0);
    signal send_to_2_490 : std_logic_vector(0 downto 0);
    signal send_to_3_495 : std_logic_vector(0 downto 0);
    signal sh_start_405 : std_logic_vector(63 downto 0);
    signal start_add_451_buffered : std_logic_vector(63 downto 0);
    signal start_next_445 : std_logic_vector(7 downto 0);
    signal type_cast_420_wire : std_logic_vector(63 downto 0);
    signal type_cast_428_wire : std_logic_vector(63 downto 0);
    signal type_cast_434_wire : std_logic_vector(63 downto 0);
    signal var_val_477 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_410_constant_part_of_offset <= "00000000000000";
    array_obj_ref_410_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_410_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_410_resized_base_address <= "00000000000000";
    array_obj_ref_521_constant_part_of_offset <= "00000000000000";
    array_obj_ref_521_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_521_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_521_resized_base_address <= "00000000000000";
    konst_397_wire_constant <= "0000000000000001";
    konst_403_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_426_wire_constant <= "0000000000000001";
    konst_439_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_459_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_461_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_469_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_510_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_519_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_547_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_415_word_offset_0 <= "00000000000000";
    ptr_deref_530_word_offset_0 <= "00000000000000";
    phi_stmt_449: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= start_add_451_buffered & nmycount_471_452_buffered;
      req <= phi_stmt_449_req_0 & phi_stmt_449_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_449",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_449_ack_0,
          idata => idata,
          odata => mycount_449,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_449
    phi_stmt_453: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_543_455_buffered & my_fetch_416_456_buffered;
      req <= phi_stmt_453_req_0 & phi_stmt_453_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_453",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_453_ack_0,
          idata => idata,
          odata => fetch_val_453,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_453
    -- flow-through select operator MUX_542_inst
    nfetch_val_543 <= fv_531 when (fn_494_delayed_13_0_534(0) /=  '0') else fetch_val_496_delayed_13_0_537;
    W_fetch_val_496_delayed_13_0_535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_496_delayed_13_0_535_inst_req_0;
      W_fetch_val_496_delayed_13_0_535_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_496_delayed_13_0_535_inst_req_1;
      W_fetch_val_496_delayed_13_0_535_inst_ack_1<= rack(0);
      W_fetch_val_496_delayed_13_0_535_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_496_delayed_13_0_535_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_496_delayed_13_0_537,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_488_delayed_7_0_524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_488_delayed_7_0_524_inst_req_0;
      W_fn_488_delayed_7_0_524_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_488_delayed_7_0_524_inst_req_1;
      W_fn_488_delayed_7_0_524_inst_ack_1<= rack(0);
      W_fn_488_delayed_7_0_524_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_488_delayed_7_0_524_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_514,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_488_delayed_7_0_526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_494_delayed_13_0_532_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_494_delayed_13_0_532_inst_req_0;
      W_fn_494_delayed_13_0_532_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_494_delayed_13_0_532_inst_req_1;
      W_fn_494_delayed_13_0_532_inst_ack_1<= rack(0);
      W_fn_494_delayed_13_0_532_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_494_delayed_13_0_532_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_514,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_494_delayed_13_0_534,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_411_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_411_final_reg_req_0;
      addr_of_411_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_411_final_reg_req_1;
      addr_of_411_final_reg_ack_1<= rack(0);
      addr_of_411_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_411_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_410_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_522_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_522_final_reg_req_0;
      addr_of_522_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_522_final_reg_req_1;
      addr_of_522_final_reg_ack_1<= rack(0);
      addr_of_522_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_522_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_521_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_416_456_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_416_456_buf_req_0;
      my_fetch_416_456_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_416_456_buf_req_1;
      my_fetch_416_456_buf_ack_1<= rack(0);
      my_fetch_416_456_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_416_456_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_416_456_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_543_455_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_543_455_buf_req_0;
      nfetch_val_543_455_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_543_455_buf_req_1;
      nfetch_val_543_455_buf_ack_1<= rack(0);
      nfetch_val_543_455_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_543_455_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_543,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_543_455_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_471_452_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_471_452_buf_req_0;
      nmycount_471_452_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_471_452_buf_req_1;
      nmycount_471_452_buf_ack_1<= rack(0);
      nmycount_471_452_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_471_452_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_471,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_471_452_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_451_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_451_buf_req_0;
      start_add_451_buf_ack_0<= wack(0);
      rreq(0) <= start_add_451_buf_req_1;
      start_add_451_buf_ack_1<= rack(0);
      start_add_451_buf : InterlockBuffer generic map ( -- 
        name => "start_add_451_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_451_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_420_inst
    process(row_size_400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_400(15 downto 0);
      type_cast_420_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_428_inst
    process(SHL_u16_u16_427_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := SHL_u16_u16_427_wire(15 downto 0);
      type_cast_428_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_434_inst
    process(row_size_400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_400(15 downto 0);
      type_cast_434_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_476_inst
    process(LSHR_u64_u64_475_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_475_wire(15 downto 0);
      var_val_477 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_410_index_1_rename
    process(R_sh_start_409_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_409_resized;
      ov(13 downto 0) := iv;
      R_sh_start_409_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_410_index_1_resize
    process(sh_start_405) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_405;
      ov := iv(13 downto 0);
      R_sh_start_409_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_410_root_address_inst
    process(array_obj_ref_410_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_410_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_410_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_521_index_1_rename
    process(LSHR_u64_u64_520_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_520_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_520_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_521_index_1_resize
    process(LSHR_u64_u64_520_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_520_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_520_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_521_root_address_inst
    process(array_obj_ref_521_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_521_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_521_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_415_addr_0
    process(ptr_deref_415_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_415_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_415_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_415_base_resize
    process(fetch_addr_412) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_412;
      ov := iv(13 downto 0);
      ptr_deref_415_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_415_gather_scatter
    process(ptr_deref_415_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_415_data_0;
      ov(63 downto 0) := iv;
      my_fetch_416 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_415_root_address_inst
    process(ptr_deref_415_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_415_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_415_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_530_addr_0
    process(ptr_deref_530_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_530_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_530_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_530_base_resize
    process(fetch_addr_523) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_523;
      ov := iv(13 downto 0);
      ptr_deref_530_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_530_gather_scatter
    process(ptr_deref_530_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_530_data_0;
      ov(63 downto 0) := iv;
      fv_531 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_530_root_address_inst
    process(ptr_deref_530_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_530_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_530_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_447_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_549_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_447_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_447_branch_req_0,
          ack0 => do_while_stmt_447_branch_ack_0,
          ack1 => do_while_stmt_447_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_399_inst
    process(num_chl_buffer, SHL_u16_u16_398_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_chl_buffer, SHL_u16_u16_398_wire, tmp_var);
      row_size_400 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_421_inst
    process(start_add_buffer, type_cast_420_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_420_wire, tmp_var);
      ea1_422 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_429_inst
    process(start_add_buffer, type_cast_428_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_428_wire, tmp_var);
      ea2_430 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_435_inst
    process(ea2_430, type_cast_434_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ea2_430, type_cast_434_wire, tmp_var);
      ea3_436 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_470_inst
    process(mycount_449) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_449, konst_469_wire_constant, tmp_var);
      nmycount_471 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_489_inst
    process(NOT_u1_u1_485_wire, ULT_u64_u1_488_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_485_wire, ULT_u64_u1_488_wire, tmp_var);
      send_to_2_490 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_462_inst
    process(mycount_449) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_449, konst_461_wire_constant, tmp_var);
      AND_u64_u64_462_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_511_inst
    process(nmycount_471) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_471, konst_510_wire_constant, tmp_var);
      AND_u64_u64_511_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_440_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_439_wire_constant, tmp_var);
      first_fill_441 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_513_inst
    process(AND_u64_u64_511_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_511_wire, konst_512_wire_constant, tmp_var);
      fn_514 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_404_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_403_wire_constant, tmp_var);
      sh_start_405 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_475_inst
    process(fetch_val_453, my_num1_466) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_453, my_num1_466, tmp_var);
      LSHR_u64_u64_475_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_520_inst
    process(nmycount_471) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_471, konst_519_wire_constant, tmp_var);
      LSHR_u64_u64_520_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_485_inst
    process(send_to_1_482) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", send_to_1_482, tmp_var);
      NOT_u1_u1_485_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u16_u16_398_inst
    process(num_chl_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(num_chl_buffer, konst_397_wire_constant, tmp_var);
      SHL_u16_u16_398_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_427_inst
    process(row_size_400) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(row_size_400, konst_426_wire_constant, tmp_var);
      SHL_u16_u16_427_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_465_inst
    process(SUB_u64_u64_463_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_463_wire, konst_464_wire_constant, tmp_var);
      my_num1_466 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_463_inst
    process(konst_459_wire_constant, AND_u64_u64_462_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_459_wire_constant, AND_u64_u64_462_wire, tmp_var);
      SUB_u64_u64_463_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_548_inst
    process(ea3_436) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(ea3_436, konst_547_wire_constant, tmp_var);
      SUB_u64_u64_548_wire <= tmp_var; --
    end process;
    -- binary operator UGE_u64_u1_494_inst
    process(mycount_449, ea2_430) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(mycount_449, ea2_430, tmp_var);
      send_to_3_495 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_481_inst
    process(mycount_449, ea1_422) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_449, ea1_422, tmp_var);
      send_to_1_482 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_488_inst
    process(mycount_449, ea2_430) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_449, ea2_430, tmp_var);
      ULT_u64_u1_488_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_549_inst
    process(mycount_449, SUB_u64_u64_548_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_449, SUB_u64_u64_548_wire, tmp_var);
      ULT_u64_u1_549_wire <= tmp_var; --
    end process;
    -- shared split operator group (23) : array_obj_ref_410_index_offset 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_409_scaled;
      array_obj_ref_410_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_410_index_offset_req_0;
      array_obj_ref_410_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_410_index_offset_req_1;
      array_obj_ref_410_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_23_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : array_obj_ref_521_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_520_scaled;
      array_obj_ref_521_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_521_index_offset_req_0;
      array_obj_ref_521_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_521_index_offset_req_1;
      array_obj_ref_521_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : ptr_deref_530_load_0 ptr_deref_415_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_530_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_415_load_0_req_0;
      ptr_deref_530_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_415_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_530_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_415_load_0_req_1;
      ptr_deref_530_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_415_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= fn_488_delayed_7_0_526(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_530_word_address_0 & ptr_deref_415_word_address_0;
      ptr_deref_530_data_0 <= data_out(127 downto 64);
      ptr_deref_415_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_444_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_444_inst_req_0;
      RPIPE_input_done_pipe_444_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_444_inst_req_1;
      RPIPE_input_done_pipe_444_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_441(0);
      start_next_445 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_497_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_497_inst_req_0;
      WPIPE_kernel_pipe1_497_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_497_inst_req_1;
      WPIPE_kernel_pipe1_497_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_482(0);
      data_in <= var_val_477;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_501_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_501_inst_req_0;
      WPIPE_kernel_pipe2_501_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_501_inst_req_1;
      WPIPE_kernel_pipe2_501_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_490(0);
      data_in <= var_val_477;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe3_505_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe3_505_inst_req_0;
      WPIPE_kernel_pipe3_505_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe3_505_inst_req_1;
      WPIPE_kernel_pipe3_505_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_495(0);
      data_in <= var_val_477;
      kernel_pipe3_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe3_pipe_write_req(0),
          oack => kernel_pipe3_pipe_write_ack(0),
          odata => kernel_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_size_pipe_551_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_551_inst_req_0;
      WPIPE_size_pipe_551_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_551_inst_req_1;
      WPIPE_size_pipe_551_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= num_chl_buffer;
      size_pipe_write_3_gI: SplitGuardInterface generic map(name => "size_pipe_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(63 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_1767_start: Boolean;
  signal sendB_CP_1767_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_616_index_offset_ack_0 : boolean;
  signal if_stmt_570_branch_req_0 : boolean;
  signal ptr_deref_866_store_0_req_0 : boolean;
  signal addr_of_617_final_reg_req_0 : boolean;
  signal ptr_deref_887_store_0_req_0 : boolean;
  signal array_obj_ref_1008_final_reg_ack_0 : boolean;
  signal addr_of_617_final_reg_ack_0 : boolean;
  signal type_cast_625_inst_req_0 : boolean;
  signal type_cast_635_inst_ack_0 : boolean;
  signal ptr_deref_887_store_0_ack_0 : boolean;
  signal type_cast_625_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1014_inst_req_1 : boolean;
  signal array_obj_ref_1008_index_offset_ack_0 : boolean;
  signal type_cast_675_inst_req_1 : boolean;
  signal type_cast_675_inst_ack_1 : boolean;
  signal ptr_deref_866_store_0_ack_1 : boolean;
  signal ptr_deref_1012_load_0_ack_0 : boolean;
  signal type_cast_645_inst_req_0 : boolean;
  signal array_obj_ref_1008_index_offset_req_1 : boolean;
  signal array_obj_ref_996_index_offset_req_1 : boolean;
  signal type_cast_675_inst_req_0 : boolean;
  signal type_cast_675_inst_ack_0 : boolean;
  signal ptr_deref_866_store_0_ack_0 : boolean;
  signal type_cast_645_inst_ack_0 : boolean;
  signal ptr_deref_887_store_0_req_1 : boolean;
  signal array_obj_ref_1008_index_offset_ack_1 : boolean;
  signal type_cast_665_inst_req_1 : boolean;
  signal type_cast_625_inst_ack_1 : boolean;
  signal type_cast_625_inst_ack_0 : boolean;
  signal type_cast_665_inst_req_0 : boolean;
  signal type_cast_665_inst_ack_0 : boolean;
  signal type_cast_665_inst_ack_1 : boolean;
  signal type_cast_856_inst_req_0 : boolean;
  signal if_stmt_570_branch_ack_1 : boolean;
  signal type_cast_635_inst_req_1 : boolean;
  signal array_obj_ref_616_index_offset_req_0 : boolean;
  signal type_cast_856_inst_ack_1 : boolean;
  signal array_obj_ref_616_index_offset_ack_1 : boolean;
  signal array_obj_ref_616_index_offset_req_1 : boolean;
  signal array_obj_ref_996_index_offset_ack_1 : boolean;
  signal type_cast_856_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1014_inst_ack_1 : boolean;
  signal type_cast_645_inst_ack_1 : boolean;
  signal type_cast_645_inst_req_1 : boolean;
  signal ptr_deref_887_store_0_ack_1 : boolean;
  signal type_cast_856_inst_req_1 : boolean;
  signal if_stmt_570_branch_ack_0 : boolean;
  signal type_cast_655_inst_req_0 : boolean;
  signal type_cast_655_inst_ack_1 : boolean;
  signal type_cast_655_inst_req_1 : boolean;
  signal type_cast_655_inst_ack_0 : boolean;
  signal type_cast_635_inst_req_0 : boolean;
  signal type_cast_635_inst_ack_1 : boolean;
  signal addr_of_617_final_reg_ack_1 : boolean;
  signal ptr_deref_621_load_0_ack_1 : boolean;
  signal ptr_deref_621_load_0_req_1 : boolean;
  signal ptr_deref_621_load_0_ack_0 : boolean;
  signal ptr_deref_621_load_0_req_0 : boolean;
  signal addr_of_617_final_reg_req_1 : boolean;
  signal array_obj_ref_1008_final_reg_req_0 : boolean;
  signal if_stmt_938_branch_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1014_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1014_inst_ack_0 : boolean;
  signal if_stmt_938_branch_ack_1 : boolean;
  signal if_stmt_938_branch_ack_0 : boolean;
  signal array_obj_ref_1008_index_offset_req_0 : boolean;
  signal type_cast_685_inst_req_0 : boolean;
  signal type_cast_685_inst_ack_0 : boolean;
  signal type_cast_685_inst_req_1 : boolean;
  signal type_cast_685_inst_ack_1 : boolean;
  signal type_cast_695_inst_req_0 : boolean;
  signal type_cast_695_inst_ack_0 : boolean;
  signal type_cast_695_inst_req_1 : boolean;
  signal type_cast_695_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_697_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_697_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_697_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_697_inst_ack_1 : boolean;
  signal array_obj_ref_996_final_reg_ack_1 : boolean;
  signal ptr_deref_1012_load_0_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_700_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_700_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_700_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_700_inst_ack_1 : boolean;
  signal array_obj_ref_996_final_reg_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_703_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_703_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_703_inst_req_1 : boolean;
  signal type_cast_919_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_703_inst_ack_1 : boolean;
  signal array_obj_ref_996_index_offset_ack_0 : boolean;
  signal array_obj_ref_996_index_offset_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_706_inst_req_0 : boolean;
  signal type_cast_919_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_706_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_706_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_706_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_709_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_709_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_709_inst_req_1 : boolean;
  signal type_cast_919_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_709_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_712_inst_req_0 : boolean;
  signal type_cast_919_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_712_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_712_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_712_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_715_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_715_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_715_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_715_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_718_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_718_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_718_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_718_inst_ack_1 : boolean;
  signal if_stmt_732_branch_req_0 : boolean;
  signal ptr_deref_845_store_0_ack_1 : boolean;
  signal ptr_deref_845_store_0_req_1 : boolean;
  signal if_stmt_732_branch_ack_1 : boolean;
  signal if_stmt_732_branch_ack_0 : boolean;
  signal type_cast_898_inst_ack_1 : boolean;
  signal if_stmt_784_branch_req_0 : boolean;
  signal type_cast_898_inst_req_1 : boolean;
  signal if_stmt_784_branch_ack_1 : boolean;
  signal ptr_deref_845_store_0_ack_0 : boolean;
  signal if_stmt_784_branch_ack_0 : boolean;
  signal ptr_deref_866_store_0_req_1 : boolean;
  signal type_cast_793_inst_req_0 : boolean;
  signal type_cast_793_inst_ack_0 : boolean;
  signal type_cast_793_inst_req_1 : boolean;
  signal ptr_deref_908_store_0_ack_1 : boolean;
  signal type_cast_793_inst_ack_1 : boolean;
  signal ptr_deref_929_store_0_ack_1 : boolean;
  signal ptr_deref_929_store_0_req_1 : boolean;
  signal type_cast_898_inst_ack_0 : boolean;
  signal array_obj_ref_799_index_offset_req_0 : boolean;
  signal ptr_deref_908_store_0_req_1 : boolean;
  signal array_obj_ref_799_index_offset_ack_0 : boolean;
  signal array_obj_ref_799_index_offset_req_1 : boolean;
  signal array_obj_ref_799_index_offset_ack_1 : boolean;
  signal array_obj_ref_996_final_reg_ack_0 : boolean;
  signal array_obj_ref_1008_final_reg_ack_1 : boolean;
  signal array_obj_ref_1008_final_reg_req_1 : boolean;
  signal addr_of_800_final_reg_req_0 : boolean;
  signal addr_of_800_final_reg_ack_0 : boolean;
  signal type_cast_898_inst_req_0 : boolean;
  signal addr_of_800_final_reg_req_1 : boolean;
  signal addr_of_800_final_reg_ack_1 : boolean;
  signal ptr_deref_1012_load_0_ack_1 : boolean;
  signal ptr_deref_1012_load_0_req_1 : boolean;
  signal ptr_deref_929_store_0_ack_0 : boolean;
  signal ptr_deref_929_store_0_req_0 : boolean;
  signal ptr_deref_908_store_0_ack_0 : boolean;
  signal ptr_deref_908_store_0_req_0 : boolean;
  signal ptr_deref_804_load_0_req_0 : boolean;
  signal ptr_deref_804_load_0_ack_0 : boolean;
  signal ptr_deref_845_store_0_req_0 : boolean;
  signal ptr_deref_804_load_0_req_1 : boolean;
  signal ptr_deref_804_load_0_ack_1 : boolean;
  signal array_obj_ref_996_final_reg_req_0 : boolean;
  signal type_cast_814_inst_req_0 : boolean;
  signal type_cast_814_inst_ack_0 : boolean;
  signal type_cast_814_inst_req_1 : boolean;
  signal type_cast_814_inst_ack_1 : boolean;
  signal type_cast_877_inst_ack_1 : boolean;
  signal type_cast_877_inst_req_1 : boolean;
  signal type_cast_877_inst_ack_0 : boolean;
  signal type_cast_877_inst_req_0 : boolean;
  signal ptr_deref_824_store_0_req_0 : boolean;
  signal ptr_deref_824_store_0_ack_0 : boolean;
  signal ptr_deref_824_store_0_req_1 : boolean;
  signal ptr_deref_824_store_0_ack_1 : boolean;
  signal type_cast_835_inst_req_0 : boolean;
  signal type_cast_835_inst_ack_0 : boolean;
  signal type_cast_835_inst_req_1 : boolean;
  signal type_cast_835_inst_ack_1 : boolean;
  signal ptr_deref_1019_load_0_req_0 : boolean;
  signal ptr_deref_1019_load_0_ack_0 : boolean;
  signal ptr_deref_1019_load_0_req_1 : boolean;
  signal ptr_deref_1019_load_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1021_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1021_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1021_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1021_inst_ack_1 : boolean;
  signal if_stmt_1035_branch_req_0 : boolean;
  signal if_stmt_1035_branch_ack_1 : boolean;
  signal if_stmt_1035_branch_ack_0 : boolean;
  signal phi_stmt_604_req_0 : boolean;
  signal type_cast_610_inst_req_0 : boolean;
  signal type_cast_610_inst_ack_0 : boolean;
  signal type_cast_610_inst_req_1 : boolean;
  signal type_cast_610_inst_ack_1 : boolean;
  signal phi_stmt_604_req_1 : boolean;
  signal phi_stmt_604_ack_0 : boolean;
  signal phi_stmt_764_req_0 : boolean;
  signal type_cast_770_inst_req_0 : boolean;
  signal type_cast_770_inst_ack_0 : boolean;
  signal type_cast_770_inst_req_1 : boolean;
  signal type_cast_770_inst_ack_1 : boolean;
  signal phi_stmt_764_req_1 : boolean;
  signal phi_stmt_764_ack_0 : boolean;
  signal phi_stmt_978_req_0 : boolean;
  signal type_cast_984_inst_req_0 : boolean;
  signal type_cast_984_inst_ack_0 : boolean;
  signal type_cast_984_inst_req_1 : boolean;
  signal type_cast_984_inst_ack_1 : boolean;
  signal phi_stmt_978_req_1 : boolean;
  signal phi_stmt_978_ack_0 : boolean;
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= size;
  size_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_1767_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_1767_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_1767_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_1767_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_1767: Block -- control-path 
    signal sendB_CP_1767_elements: BooleanArray(137 downto 0);
    -- 
  begin -- 
    sendB_CP_1767_elements(0) <= sendB_CP_1767_start;
    sendB_CP_1767_symbol <= sendB_CP_1767_elements(137);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_557/assign_stmt_563_to_assign_stmt_569__entry__
      -- CP-element group 0: 	 branch_block_stmt_557/if_stmt_570_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_557/assign_stmt_563_to_assign_stmt_569__exit__
      -- CP-element group 0: 	 branch_block_stmt_557/if_stmt_570_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_557/R_cmp77_571_place
      -- CP-element group 0: 	 branch_block_stmt_557/if_stmt_570__entry__
      -- CP-element group 0: 	 branch_block_stmt_557/if_stmt_570_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_557/branch_block_stmt_557__entry__
      -- CP-element group 0: 	 branch_block_stmt_557/if_stmt_570_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_557/if_stmt_570_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_557/$entry
      -- CP-element group 0: 	 branch_block_stmt_557/assign_stmt_563_to_assign_stmt_569/$exit
      -- CP-element group 0: 	 branch_block_stmt_557/assign_stmt_563_to_assign_stmt_569/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_557/if_stmt_570_else_link/$entry
      -- 
    branch_req_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(0), ack => if_stmt_570_branch_req_0); -- 
    -- CP-element group 1:  merge  transition  place  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	119 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_557/bbx_xnph_forx_xbody
      -- CP-element group 1: 	 branch_block_stmt_557/if_stmt_570_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_557/assign_stmt_582_to_assign_stmt_601/$exit
      -- CP-element group 1: 	 branch_block_stmt_557/if_stmt_570_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_557/assign_stmt_582_to_assign_stmt_601__exit__
      -- CP-element group 1: 	 branch_block_stmt_557/assign_stmt_582_to_assign_stmt_601__entry__
      -- CP-element group 1: 	 branch_block_stmt_557/assign_stmt_582_to_assign_stmt_601/$entry
      -- CP-element group 1: 	 branch_block_stmt_557/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_557/merge_stmt_576__exit__
      -- CP-element group 1: 	 branch_block_stmt_557/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_557/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_557/merge_stmt_576_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_557/merge_stmt_576_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_557/merge_stmt_576_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_557/merge_stmt_576_PhiAck/dummy
      -- CP-element group 1: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/phi_stmt_604/$entry
      -- CP-element group 1: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/$entry
      -- 
    if_choice_transition_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_570_branch_ack_1, ack => sendB_CP_1767_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	125 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_557/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_557/if_stmt_570_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_557/if_stmt_570_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/phi_stmt_764/$entry
      -- CP-element group 2: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/$entry
      -- 
    else_choice_transition_1840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_570_branch_ack_0, ack => sendB_CP_1767_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	124 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	48 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_sample_complete
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_616_index_offset_ack_0, ack => sendB_CP_1767_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	124 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (11) 
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_base_plus_offset/$entry
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_root_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_request/$entry
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_offset_calculated
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_request/req
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Update/ack
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_base_plus_offset/$exit
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_616_index_offset_ack_1, ack => sendB_CP_1767_elements(4)); -- 
    req_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(4), ack => addr_of_617_final_reg_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_request/$exit
      -- CP-element group 5: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_request/ack
      -- 
    ack_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_617_final_reg_ack_0, ack => sendB_CP_1767_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	124 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (24) 
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_word_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_address_resized
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_addr_resize/$entry
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_addr_resize/$exit
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_addr_resize/base_resize_req
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_addr_resize/base_resize_ack
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_complete/ack
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/word_access_start/word_0/rr
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/word_access_start/$entry
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_word_addrgen/root_register_ack
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_word_addrgen/root_register_req
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_word_addrgen/$exit
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_word_addrgen/$entry
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_617_final_reg_ack_1, ack => sendB_CP_1767_elements(6)); -- 
    rr_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(6), ack => ptr_deref_621_load_0_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Sample/$exit
      -- 
    ra_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_0_ack_0, ack => sendB_CP_1767_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	124 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	13 
    -- CP-element group 8: 	15 
    -- CP-element group 8: 	17 
    -- CP-element group 8: 	19 
    -- CP-element group 8:  members (33) 
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/ptr_deref_621_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/ptr_deref_621_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/ptr_deref_621_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/ptr_deref_621_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Sample/rr
      -- 
    ca_1939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_0_ack_1, ack => sendB_CP_1767_elements(8)); -- 
    rr_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_695_inst_req_0); -- 
    rr_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_625_inst_req_0); -- 
    rr_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_635_inst_req_0); -- 
    rr_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_645_inst_req_0); -- 
    rr_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_655_inst_req_0); -- 
    rr_2008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_665_inst_req_0); -- 
    rr_2022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_675_inst_req_0); -- 
    rr_2036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(8), ack => type_cast_685_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_sample_completed_
      -- 
    ra_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_625_inst_ack_0, ack => sendB_CP_1767_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	124 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	45 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_update_completed_
      -- 
    ca_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_625_inst_ack_1, ack => sendB_CP_1767_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_sample_completed_
      -- 
    ra_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_0, ack => sendB_CP_1767_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	124 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	42 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_update_completed_
      -- 
    ca_1972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_1, ack => sendB_CP_1767_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Sample/$exit
      -- 
    ra_1981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_0, ack => sendB_CP_1767_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	124 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	39 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_update_completed_
      -- 
    ca_1986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_1, ack => sendB_CP_1767_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	8 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Sample/ra
      -- 
    ra_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_655_inst_ack_0, ack => sendB_CP_1767_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	124 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	36 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Update/$exit
      -- 
    ca_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_655_inst_ack_1, ack => sendB_CP_1767_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	8 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Sample/$exit
      -- 
    ra_2009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_0, ack => sendB_CP_1767_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	124 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_update_completed_
      -- 
    ca_2014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_1, ack => sendB_CP_1767_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	8 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Sample/ra
      -- 
    ra_2023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_675_inst_ack_0, ack => sendB_CP_1767_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	124 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	30 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_update_completed_
      -- 
    ca_2028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_675_inst_ack_1, ack => sendB_CP_1767_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Sample/ra
      -- 
    ra_2037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_685_inst_ack_0, ack => sendB_CP_1767_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	124 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Update/ca
      -- 
    ca_2042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_685_inst_ack_1, ack => sendB_CP_1767_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Sample/ra
      -- 
    ra_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_0, ack => sendB_CP_1767_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	124 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Sample/req
      -- 
    ca_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_1, ack => sendB_CP_1767_elements(24)); -- 
    req_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(24), ack => WPIPE_maxpool_output_pipe_697_inst_req_0); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_update_start_
      -- CP-element group 25: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Sample/ack
      -- CP-element group 25: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Update/req
      -- 
    ack_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_697_inst_ack_0, ack => sendB_CP_1767_elements(25)); -- 
    req_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(25), ack => WPIPE_maxpool_output_pipe_697_inst_req_1); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_697_Update/ack
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_697_inst_ack_1, ack => sendB_CP_1767_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Sample/req
      -- 
    req_2078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(27), ack => WPIPE_maxpool_output_pipe_700_inst_req_0); -- 
    sendB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(22) & sendB_CP_1767_elements(26);
      gj_sendB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_update_start_
      -- CP-element group 28: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Update/req
      -- 
    ack_2079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_700_inst_ack_0, ack => sendB_CP_1767_elements(28)); -- 
    req_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(28), ack => WPIPE_maxpool_output_pipe_700_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_700_Update/ack
      -- 
    ack_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_700_inst_ack_1, ack => sendB_CP_1767_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: 	20 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Sample/req
      -- 
    req_2092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(30), ack => WPIPE_maxpool_output_pipe_703_inst_req_0); -- 
    sendB_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(29) & sendB_CP_1767_elements(20);
      gj_sendB_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_update_start_
      -- CP-element group 31: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Update/req
      -- 
    ack_2093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_703_inst_ack_0, ack => sendB_CP_1767_elements(31)); -- 
    req_2097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(31), ack => WPIPE_maxpool_output_pipe_703_inst_req_1); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_703_Update/ack
      -- 
    ack_2098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_703_inst_ack_1, ack => sendB_CP_1767_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	18 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Sample/req
      -- 
    req_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(33), ack => WPIPE_maxpool_output_pipe_706_inst_req_0); -- 
    sendB_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(32) & sendB_CP_1767_elements(18);
      gj_sendB_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_update_start_
      -- CP-element group 34: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Update/req
      -- 
    ack_2107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_706_inst_ack_0, ack => sendB_CP_1767_elements(34)); -- 
    req_2111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(34), ack => WPIPE_maxpool_output_pipe_706_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_706_Update/ack
      -- 
    ack_2112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_706_inst_ack_1, ack => sendB_CP_1767_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	16 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Sample/req
      -- 
    req_2120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(36), ack => WPIPE_maxpool_output_pipe_709_inst_req_0); -- 
    sendB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(35) & sendB_CP_1767_elements(16);
      gj_sendB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_update_start_
      -- CP-element group 37: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Update/req
      -- 
    ack_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_709_inst_ack_0, ack => sendB_CP_1767_elements(37)); -- 
    req_2125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(37), ack => WPIPE_maxpool_output_pipe_709_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_709_Update/ack
      -- 
    ack_2126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_709_inst_ack_1, ack => sendB_CP_1767_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Sample/req
      -- 
    req_2134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(39), ack => WPIPE_maxpool_output_pipe_712_inst_req_0); -- 
    sendB_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(38) & sendB_CP_1767_elements(14);
      gj_sendB_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_update_start_
      -- CP-element group 40: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Update/req
      -- 
    ack_2135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_712_inst_ack_0, ack => sendB_CP_1767_elements(40)); -- 
    req_2139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(40), ack => WPIPE_maxpool_output_pipe_712_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_712_Update/ack
      -- 
    ack_2140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_712_inst_ack_1, ack => sendB_CP_1767_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	12 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Sample/req
      -- 
    req_2148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(42), ack => WPIPE_maxpool_output_pipe_715_inst_req_0); -- 
    sendB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(41) & sendB_CP_1767_elements(12);
      gj_sendB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_update_start_
      -- CP-element group 43: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Update/req
      -- 
    ack_2149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_715_inst_ack_0, ack => sendB_CP_1767_elements(43)); -- 
    req_2153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(43), ack => WPIPE_maxpool_output_pipe_715_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_715_Update/ack
      -- 
    ack_2154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_715_inst_ack_1, ack => sendB_CP_1767_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Sample/req
      -- 
    req_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(45), ack => WPIPE_maxpool_output_pipe_718_inst_req_0); -- 
    sendB_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(44) & sendB_CP_1767_elements(10);
      gj_sendB_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_update_start_
      -- CP-element group 46: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Update/req
      -- 
    ack_2163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_718_inst_ack_0, ack => sendB_CP_1767_elements(46)); -- 
    req_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(46), ack => WPIPE_maxpool_output_pipe_718_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/WPIPE_maxpool_output_pipe_718_Update/ack
      -- 
    ack_2168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_718_inst_ack_1, ack => sendB_CP_1767_elements(47)); -- 
    -- CP-element group 48:  branch  join  transition  place  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	3 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (10) 
      -- CP-element group 48: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731__exit__
      -- CP-element group 48: 	 branch_block_stmt_557/if_stmt_732__entry__
      -- CP-element group 48: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/$exit
      -- CP-element group 48: 	 branch_block_stmt_557/if_stmt_732_dead_link/$entry
      -- CP-element group 48: 	 branch_block_stmt_557/if_stmt_732_eval_test/$entry
      -- CP-element group 48: 	 branch_block_stmt_557/if_stmt_732_eval_test/$exit
      -- CP-element group 48: 	 branch_block_stmt_557/if_stmt_732_eval_test/branch_req
      -- CP-element group 48: 	 branch_block_stmt_557/R_exitcond_733_place
      -- CP-element group 48: 	 branch_block_stmt_557/if_stmt_732_if_link/$entry
      -- CP-element group 48: 	 branch_block_stmt_557/if_stmt_732_else_link/$entry
      -- 
    branch_req_2176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(48), ack => if_stmt_732_branch_req_0); -- 
    sendB_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(47) & sendB_CP_1767_elements(3);
      gj_sendB_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	127 
    -- CP-element group 49: 	126 
    -- CP-element group 49:  members (24) 
      -- CP-element group 49: 	 branch_block_stmt_557/merge_stmt_738__exit__
      -- CP-element group 49: 	 branch_block_stmt_557/assign_stmt_745_to_assign_stmt_761__entry__
      -- CP-element group 49: 	 branch_block_stmt_557/assign_stmt_745_to_assign_stmt_761__exit__
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 49: 	 branch_block_stmt_557/if_stmt_732_if_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_557/if_stmt_732_if_link/if_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 49: 	 branch_block_stmt_557/assign_stmt_745_to_assign_stmt_761/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/assign_stmt_745_to_assign_stmt_761/$exit
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_557/merge_stmt_738_PhiReqMerge
      -- CP-element group 49: 	 branch_block_stmt_557/merge_stmt_738_PhiAck/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/merge_stmt_738_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_557/merge_stmt_738_PhiAck/dummy
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_732_branch_ack_1, ack => sendB_CP_1767_elements(49)); -- 
    rr_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(49), ack => type_cast_770_inst_req_0); -- 
    cr_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(49), ack => type_cast_770_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  place  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	120 
    -- CP-element group 50: 	121 
    -- CP-element group 50:  members (12) 
      -- CP-element group 50: 	 branch_block_stmt_557/if_stmt_732_else_link/$exit
      -- CP-element group 50: 	 branch_block_stmt_557/if_stmt_732_else_link/else_choice_transition
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/$entry
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/$entry
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/$entry
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/$entry
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_732_branch_ack_0, ack => sendB_CP_1767_elements(50)); -- 
    rr_3022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(50), ack => type_cast_610_inst_req_0); -- 
    cr_3027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(50), ack => type_cast_610_inst_req_1); -- 
    -- CP-element group 51:  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	130 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	137 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_557/if_stmt_784_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_557/if_stmt_784_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_557/forx_xend_sendRemainingElementsx_xexit
      -- CP-element group 51: 	 branch_block_stmt_557/forx_xend_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_557/forx_xend_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_784_branch_ack_1, ack => sendB_CP_1767_elements(51)); -- 
    -- CP-element group 52:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	130 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	80 
    -- CP-element group 52: 	88 
    -- CP-element group 52: 	82 
    -- CP-element group 52: 	83 
    -- CP-element group 52: 	87 
    -- CP-element group 52: 	65 
    -- CP-element group 52: 	67 
    -- CP-element group 52: 	85 
    -- CP-element group 52: 	60 
    -- CP-element group 52: 	62 
    -- CP-element group 52: 	63 
    -- CP-element group 52: 	90 
    -- CP-element group 52: 	68 
    -- CP-element group 52: 	70 
    -- CP-element group 52: 	72 
    -- CP-element group 52: 	73 
    -- CP-element group 52: 	75 
    -- CP-element group 52: 	77 
    -- CP-element group 52: 	78 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52: 	56 
    -- CP-element group 52: 	58 
    -- CP-element group 52:  members (186) 
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937__entry__
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/merge_stmt_790__exit__
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/if_stmt_784_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/if_stmt_784_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_557/forx_xend_ifx_xthen
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_resized_1
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_scaled_1
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_computed_1
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_resize_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_resize_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_resize_1/index_resize_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_resize_1/index_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_scale_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_scale_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_scale_1/scale_rename_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_index_scale_1/scale_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_update_start
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Update/req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_complete/req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_update_start_
      -- CP-element group 52: 	 branch_block_stmt_557/forx_xend_ifx_xthen_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/forx_xend_ifx_xthen_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/merge_stmt_790_PhiReqMerge
      -- CP-element group 52: 	 branch_block_stmt_557/merge_stmt_790_PhiAck/$entry
      -- CP-element group 52: 	 branch_block_stmt_557/merge_stmt_790_PhiAck/$exit
      -- CP-element group 52: 	 branch_block_stmt_557/merge_stmt_790_PhiAck/dummy
      -- 
    else_choice_transition_2210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_784_branch_ack_0, ack => sendB_CP_1767_elements(52)); -- 
    cr_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => ptr_deref_887_store_0_req_1); -- 
    cr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_856_inst_req_1); -- 
    cr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_919_inst_req_1); -- 
    cr_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => ptr_deref_845_store_0_req_1); -- 
    cr_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_898_inst_req_1); -- 
    cr_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => ptr_deref_866_store_0_req_1); -- 
    rr_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_793_inst_req_0); -- 
    cr_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_793_inst_req_1); -- 
    cr_2708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => ptr_deref_929_store_0_req_1); -- 
    req_2254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => array_obj_ref_799_index_offset_req_0); -- 
    cr_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => ptr_deref_908_store_0_req_1); -- 
    req_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => array_obj_ref_799_index_offset_req_1); -- 
    req_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => addr_of_800_final_reg_req_1); -- 
    cr_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => ptr_deref_804_load_0_req_1); -- 
    cr_2338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_814_inst_req_1); -- 
    cr_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_877_inst_req_1); -- 
    cr_2388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => ptr_deref_824_store_0_req_1); -- 
    cr_2402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(52), ack => type_cast_835_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Sample/ra
      -- 
    ra_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_0, ack => sendB_CP_1767_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	96 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_793_Update/ca
      -- 
    ca_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_1, ack => sendB_CP_1767_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	96 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_sample_complete
      -- CP-element group 55: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Sample/ack
      -- 
    ack_2255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_799_index_offset_ack_0, ack => sendB_CP_1767_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (11) 
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_offset_calculated
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_final_index_sum_regn_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/array_obj_ref_799_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_request/$entry
      -- CP-element group 56: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_request/req
      -- 
    ack_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_799_index_offset_ack_1, ack => sendB_CP_1767_elements(56)); -- 
    req_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(56), ack => addr_of_800_final_reg_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_request/$exit
      -- CP-element group 57: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_request/ack
      -- 
    ack_2270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_800_final_reg_ack_0, ack => sendB_CP_1767_elements(57)); -- 
    -- CP-element group 58:  join  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	52 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_complete/$exit
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/addr_of_800_complete/ack
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/word_access_start/word_0/rr
      -- 
    ack_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_800_final_reg_ack_1, ack => sendB_CP_1767_elements(58)); -- 
    rr_2308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(58), ack => ptr_deref_804_load_0_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Sample/word_access_start/word_0/ra
      -- 
    ra_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_804_load_0_ack_0, ack => sendB_CP_1767_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	52 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	81 
    -- CP-element group 60: 	86 
    -- CP-element group 60: 	66 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	71 
    -- CP-element group 60: 	76 
    -- CP-element group 60:  members (27) 
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/ptr_deref_804_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/ptr_deref_804_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/ptr_deref_804_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_804_Update/ptr_deref_804_Merge/merge_ack
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Sample/rr
      -- 
    ca_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_804_load_0_ack_1, ack => sendB_CP_1767_elements(60)); -- 
    rr_2589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(60), ack => type_cast_898_inst_req_0); -- 
    rr_2397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(60), ack => type_cast_835_inst_req_0); -- 
    rr_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(60), ack => type_cast_814_inst_req_0); -- 
    rr_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(60), ack => type_cast_919_inst_req_0); -- 
    rr_2461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(60), ack => type_cast_856_inst_req_0); -- 
    rr_2525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(60), ack => type_cast_877_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Sample/ra
      -- 
    ra_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_0, ack => sendB_CP_1767_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	52 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_814_Update/ca
      -- 
    ca_2339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_1, ack => sendB_CP_1767_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: 	52 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/ptr_deref_824_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/ptr_deref_824_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/ptr_deref_824_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/ptr_deref_824_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/word_access_start/word_0/rr
      -- 
    rr_2377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(63), ack => ptr_deref_824_store_0_req_0); -- 
    sendB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(62) & sendB_CP_1767_elements(52);
      gj_sendB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	91 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Sample/word_access_start/word_0/ra
      -- 
    ra_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_824_store_0_ack_0, ack => sendB_CP_1767_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	52 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	96 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_Update/word_access_complete/word_0/ca
      -- 
    ca_2389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_824_store_0_ack_1, ack => sendB_CP_1767_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Sample/ra
      -- 
    ra_2398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_0, ack => sendB_CP_1767_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	52 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_835_Update/ca
      -- 
    ca_2403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_1, ack => sendB_CP_1767_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: 	91 
    -- CP-element group 68: 	52 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (9) 
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/word_access_start/word_0/$entry
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/ptr_deref_845_Split/split_req
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/ptr_deref_845_Split/$exit
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/ptr_deref_845_Split/split_ack
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/ptr_deref_845_Split/$entry
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/word_access_start/$entry
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/word_access_start/word_0/rr
      -- CP-element group 68: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_sample_start_
      -- 
    rr_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(68), ack => ptr_deref_845_store_0_req_0); -- 
    sendB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(67) & sendB_CP_1767_elements(91) & sendB_CP_1767_elements(52);
      gj_sendB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	92 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/word_access_start/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/word_access_start/$exit
      -- CP-element group 69: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Sample/word_access_start/word_0/ra
      -- CP-element group 69: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_sample_completed_
      -- 
    ra_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_845_store_0_ack_0, ack => sendB_CP_1767_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	52 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	96 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/word_access_complete/word_0/ca
      -- CP-element group 70: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/word_access_complete/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/word_access_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_update_completed_
      -- 
    ca_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_845_store_0_ack_1, ack => sendB_CP_1767_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	60 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_sample_completed_
      -- 
    ra_2462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_856_inst_ack_0, ack => sendB_CP_1767_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	52 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_856_update_completed_
      -- 
    ca_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_856_inst_ack_1, ack => sendB_CP_1767_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	92 
    -- CP-element group 73: 	72 
    -- CP-element group 73: 	52 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/ptr_deref_866_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/ptr_deref_866_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/ptr_deref_866_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/ptr_deref_866_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/$entry
      -- 
    rr_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(73), ack => ptr_deref_866_store_0_req_0); -- 
    sendB_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(92) & sendB_CP_1767_elements(72) & sendB_CP_1767_elements(52);
      gj_sendB_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	93 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/word_access_start/word_0/ra
      -- CP-element group 74: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Sample/$exit
      -- 
    ra_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_866_store_0_ack_0, ack => sendB_CP_1767_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	96 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/word_access_complete/word_0/ca
      -- CP-element group 75: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_Update/word_access_complete/$exit
      -- 
    ca_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_866_store_0_ack_1, ack => sendB_CP_1767_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	60 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Sample/ra
      -- 
    ra_2526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_877_inst_ack_0, ack => sendB_CP_1767_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	52 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_877_Update/$exit
      -- 
    ca_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_877_inst_ack_1, ack => sendB_CP_1767_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	77 
    -- CP-element group 78: 	52 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/word_access_start/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/word_access_start/word_0/rr
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/word_access_start/$entry
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/ptr_deref_887_Split/split_ack
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/ptr_deref_887_Split/split_req
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/ptr_deref_887_Split/$exit
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/ptr_deref_887_Split/$entry
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_sample_start_
      -- 
    rr_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(78), ack => ptr_deref_887_store_0_req_0); -- 
    sendB_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(93) & sendB_CP_1767_elements(77) & sendB_CP_1767_elements(52);
      gj_sendB_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	94 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/word_access_start/word_0/ra
      -- CP-element group 79: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/word_access_start/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/word_access_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_sample_completed_
      -- 
    ra_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_887_store_0_ack_0, ack => sendB_CP_1767_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	52 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	96 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/word_access_complete/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/word_access_complete/word_0/ca
      -- CP-element group 80: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_Update/word_access_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_update_completed_
      -- 
    ca_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_887_store_0_ack_1, ack => sendB_CP_1767_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	60 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Sample/$exit
      -- 
    ra_2590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_0, ack => sendB_CP_1767_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	52 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_898_Update/$exit
      -- 
    ca_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_1, ack => sendB_CP_1767_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: 	94 
    -- CP-element group 83: 	52 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/ptr_deref_908_Split/$entry
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/word_access_start/word_0/rr
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/word_access_start/word_0/$entry
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/word_access_start/$entry
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/ptr_deref_908_Split/split_ack
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/ptr_deref_908_Split/split_req
      -- CP-element group 83: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/ptr_deref_908_Split/$exit
      -- 
    rr_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(83), ack => ptr_deref_908_store_0_req_0); -- 
    sendB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(82) & sendB_CP_1767_elements(94) & sendB_CP_1767_elements(52);
      gj_sendB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	95 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/word_access_start/word_0/ra
      -- CP-element group 84: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/word_access_start/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Sample/word_access_start/$exit
      -- 
    ra_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_908_store_0_ack_0, ack => sendB_CP_1767_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	52 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	96 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/word_access_complete/word_0/ca
      -- CP-element group 85: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/word_access_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_Update/$exit
      -- 
    ca_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_908_store_0_ack_1, ack => sendB_CP_1767_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	60 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_sample_completed_
      -- 
    ra_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_919_inst_ack_0, ack => sendB_CP_1767_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	52 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/type_cast_919_update_completed_
      -- 
    ca_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_919_inst_ack_1, ack => sendB_CP_1767_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: 	95 
    -- CP-element group 88: 	52 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/ptr_deref_929_Split/$entry
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/word_access_start/word_0/rr
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/word_access_start/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/word_access_start/$entry
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/ptr_deref_929_Split/split_ack
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/ptr_deref_929_Split/split_req
      -- CP-element group 88: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/ptr_deref_929_Split/$exit
      -- 
    rr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(88), ack => ptr_deref_929_store_0_req_0); -- 
    sendB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(87) & sendB_CP_1767_elements(95) & sendB_CP_1767_elements(52);
      gj_sendB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/word_access_start/word_0/ra
      -- CP-element group 89: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/word_access_start/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Sample/word_access_start/$exit
      -- 
    ra_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_929_store_0_ack_0, ack => sendB_CP_1767_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	52 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	96 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/word_access_complete/word_0/ca
      -- CP-element group 90: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/word_access_complete/word_0/$exit
      -- CP-element group 90: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/word_access_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_929_Update/$exit
      -- 
    ca_2709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_929_store_0_ack_1, ack => sendB_CP_1767_elements(90)); -- 
    -- CP-element group 91:  transition  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	64 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	68 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_824_ptr_deref_845_delay
      -- 
    -- Element group sendB_CP_1767_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(64), ack => sendB_CP_1767_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	69 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	73 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_845_ptr_deref_866_delay
      -- 
    -- Element group sendB_CP_1767_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(69), ack => sendB_CP_1767_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  transition  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	74 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	78 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_866_ptr_deref_887_delay
      -- 
    -- Element group sendB_CP_1767_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(74), ack => sendB_CP_1767_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  transition  delay-element  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	79 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	83 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_887_ptr_deref_908_delay
      -- 
    -- Element group sendB_CP_1767_elements(94) is a control-delay.
    cp_element_94_delay: control_delay_element  generic map(name => " 94_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(79), ack => sendB_CP_1767_elements(94), clk => clk, reset =>reset);
    -- CP-element group 95:  transition  delay-element  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	84 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	88 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/ptr_deref_908_ptr_deref_929_delay
      -- 
    -- Element group sendB_CP_1767_elements(95) is a control-delay.
    cp_element_95_delay: control_delay_element  generic map(name => " 95_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(84), ack => sendB_CP_1767_elements(95), clk => clk, reset =>reset);
    -- CP-element group 96:  branch  join  transition  place  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	80 
    -- CP-element group 96: 	65 
    -- CP-element group 96: 	85 
    -- CP-element group 96: 	90 
    -- CP-element group 96: 	70 
    -- CP-element group 96: 	75 
    -- CP-element group 96: 	54 
    -- CP-element group 96: 	55 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (10) 
      -- CP-element group 96: 	 branch_block_stmt_557/if_stmt_938_dead_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_557/if_stmt_938_eval_test/$entry
      -- CP-element group 96: 	 branch_block_stmt_557/if_stmt_938__entry__
      -- CP-element group 96: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937__exit__
      -- CP-element group 96: 	 branch_block_stmt_557/if_stmt_938_else_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_557/if_stmt_938_eval_test/$exit
      -- CP-element group 96: 	 branch_block_stmt_557/if_stmt_938_eval_test/branch_req
      -- CP-element group 96: 	 branch_block_stmt_557/if_stmt_938_if_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_557/assign_stmt_794_to_assign_stmt_937/$exit
      -- CP-element group 96: 	 branch_block_stmt_557/R_cmp53x_xi_939_place
      -- 
    branch_req_2722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(96), ack => if_stmt_938_branch_req_0); -- 
    sendB_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(80) & sendB_CP_1767_elements(65) & sendB_CP_1767_elements(85) & sendB_CP_1767_elements(90) & sendB_CP_1767_elements(70) & sendB_CP_1767_elements(75) & sendB_CP_1767_elements(54) & sendB_CP_1767_elements(55);
      gj_sendB_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  place  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	137 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_557/if_stmt_938_if_link/$exit
      -- CP-element group 97: 	 branch_block_stmt_557/if_stmt_938_if_link/if_choice_transition
      -- CP-element group 97: 	 branch_block_stmt_557/ifx_xthen_sendRemainingElementsx_xexit
      -- CP-element group 97: 	 branch_block_stmt_557/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 97: 	 branch_block_stmt_557/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_938_branch_ack_1, ack => sendB_CP_1767_elements(97)); -- 
    -- CP-element group 98:  merge  transition  place  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	131 
    -- CP-element group 98:  members (18) 
      -- CP-element group 98: 	 branch_block_stmt_557/assign_stmt_950_to_assign_stmt_975/$exit
      -- CP-element group 98: 	 branch_block_stmt_557/assign_stmt_950_to_assign_stmt_975__exit__
      -- CP-element group 98: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 98: 	 branch_block_stmt_557/assign_stmt_950_to_assign_stmt_975__entry__
      -- CP-element group 98: 	 branch_block_stmt_557/merge_stmt_944__exit__
      -- CP-element group 98: 	 branch_block_stmt_557/assign_stmt_950_to_assign_stmt_975/$entry
      -- CP-element group 98: 	 branch_block_stmt_557/ifx_xthen_bbx_xnphx_xi
      -- CP-element group 98: 	 branch_block_stmt_557/if_stmt_938_else_link/$exit
      -- CP-element group 98: 	 branch_block_stmt_557/if_stmt_938_else_link/else_choice_transition
      -- CP-element group 98: 	 branch_block_stmt_557/ifx_xthen_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 98: 	 branch_block_stmt_557/ifx_xthen_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 98: 	 branch_block_stmt_557/merge_stmt_944_PhiReqMerge
      -- CP-element group 98: 	 branch_block_stmt_557/merge_stmt_944_PhiAck/$entry
      -- CP-element group 98: 	 branch_block_stmt_557/merge_stmt_944_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_557/merge_stmt_944_PhiAck/dummy
      -- CP-element group 98: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 98: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/$entry
      -- CP-element group 98: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/$entry
      -- 
    else_choice_transition_2731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_938_branch_ack_0, ack => sendB_CP_1767_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	136 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	116 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_sample_complete
      -- 
    ack_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_996_index_offset_ack_0, ack => sendB_CP_1767_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	136 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (11) 
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_request/$entry
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_base_plus_offset/$exit
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_base_plus_offset/$entry
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_base_plus_offset/sum_rename_ack
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_base_plus_offset/sum_rename_req
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_offset_calculated
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_root_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_request/req
      -- 
    ack_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_996_index_offset_ack_1, ack => sendB_CP_1767_elements(100)); -- 
    req_2780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(100), ack => array_obj_ref_996_final_reg_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_request/$exit
      -- CP-element group 101: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_request/ack
      -- 
    ack_2781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_996_final_reg_ack_0, ack => sendB_CP_1767_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	136 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	107 
    -- CP-element group 102:  members (24) 
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_complete/ack
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/word_access_start/word_0/rr
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/word_access_start/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/word_access_start/$entry
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_word_addrgen/root_register_ack
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_word_addrgen/root_register_req
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_word_addrgen/$exit
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_word_addrgen/$entry
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_plus_offset/sum_rename_ack
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_plus_offset/sum_rename_req
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_plus_offset/$exit
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_plus_offset/$entry
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_addr_resize/base_resize_ack
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_addr_resize/base_resize_req
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_addr_resize/$exit
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_addr_resize/$entry
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_address_resized
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_root_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_word_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_base_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_update_completed_
      -- 
    ack_2786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_996_final_reg_ack_1, ack => sendB_CP_1767_elements(102)); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(102), ack => ptr_deref_1012_load_0_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	136 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	116 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Sample/ack
      -- CP-element group 103: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_sample_complete
      -- 
    ack_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_index_offset_ack_0, ack => sendB_CP_1767_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	136 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (11) 
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_base_plus_offset/$entry
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_base_plus_offset/sum_rename_ack
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_base_plus_offset/sum_rename_req
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_base_plus_offset/$exit
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_request/$entry
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_request/req
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_offset_calculated
      -- CP-element group 104: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_root_address_calculated
      -- 
    ack_2818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_index_offset_ack_1, ack => sendB_CP_1767_elements(104)); -- 
    req_2827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(104), ack => array_obj_ref_1008_final_reg_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_request/ack
      -- CP-element group 105: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_request/$exit
      -- CP-element group 105: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_sample_completed_
      -- 
    ack_2828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_final_reg_ack_0, ack => sendB_CP_1767_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	136 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	111 
    -- CP-element group 106:  members (24) 
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_complete/$exit
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_word_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_word_addrgen/root_register_req
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_word_addrgen/$entry
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_addr_resize/$entry
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_word_addrgen/$exit
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_addr_resize/base_resize_ack
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_addr_resize/base_resize_req
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_addr_resize/$exit
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_address_resized
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_root_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_plus_offset/sum_rename_ack
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_complete/ack
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_plus_offset/sum_rename_req
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_plus_offset/$entry
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_base_plus_offset/$exit
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_word_addrgen/root_register_ack
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/word_access_start/$entry
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/word_access_start/word_0/$entry
      -- CP-element group 106: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/word_access_start/word_0/rr
      -- 
    ack_2833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_final_reg_ack_1, ack => sendB_CP_1767_elements(106)); -- 
    rr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(106), ack => ptr_deref_1019_load_0_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	102 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/word_access_start/word_0/ra
      -- CP-element group 107: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/word_access_start/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/word_access_start/$exit
      -- CP-element group 107: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_sample_completed_
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1012_load_0_ack_0, ack => sendB_CP_1767_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	136 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (12) 
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Sample/req
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/ptr_deref_1012_Merge/merge_ack
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/ptr_deref_1012_Merge/merge_req
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/ptr_deref_1012_Merge/$exit
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/ptr_deref_1012_Merge/$entry
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/word_access_complete/word_0/ca
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/word_access_complete/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/word_access_complete/$exit
      -- 
    ca_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1012_load_0_ack_1, ack => sendB_CP_1767_elements(108)); -- 
    req_2891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(108), ack => WPIPE_maxpool_output_pipe_1014_inst_req_0); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Update/req
      -- CP-element group 109: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_update_start_
      -- CP-element group 109: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Sample/ack
      -- CP-element group 109: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_sample_completed_
      -- 
    ack_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1014_inst_ack_0, ack => sendB_CP_1767_elements(109)); -- 
    req_2896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(109), ack => WPIPE_maxpool_output_pipe_1014_inst_req_1); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_Update/ack
      -- CP-element group 110: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1014_update_completed_
      -- 
    ack_2897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1014_inst_ack_1, ack => sendB_CP_1767_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	106 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/word_access_start/$exit
      -- CP-element group 111: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/word_access_start/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Sample/word_access_start/word_0/ra
      -- 
    ra_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1019_load_0_ack_0, ack => sendB_CP_1767_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	136 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/word_access_complete/$exit
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/word_access_complete/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/word_access_complete/word_0/ca
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/ptr_deref_1019_Merge/$entry
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/ptr_deref_1019_Merge/$exit
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/ptr_deref_1019_Merge/merge_req
      -- CP-element group 112: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/ptr_deref_1019_Merge/merge_ack
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1019_load_0_ack_1, ack => sendB_CP_1767_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Sample/req
      -- 
    req_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(113), ack => WPIPE_maxpool_output_pipe_1021_inst_req_0); -- 
    sendB_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(110) & sendB_CP_1767_elements(112);
      gj_sendB_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_update_start_
      -- CP-element group 114: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Update/req
      -- 
    ack_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1021_inst_ack_0, ack => sendB_CP_1767_elements(114)); -- 
    req_2960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(114), ack => WPIPE_maxpool_output_pipe_1021_inst_req_1); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/WPIPE_maxpool_output_pipe_1021_Update/ack
      -- 
    ack_2961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1021_inst_ack_1, ack => sendB_CP_1767_elements(115)); -- 
    -- CP-element group 116:  branch  join  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: 	103 
    -- CP-element group 116: 	99 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/$exit
      -- CP-element group 116: 	 branch_block_stmt_557/if_stmt_1035__entry__
      -- CP-element group 116: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034__exit__
      -- CP-element group 116: 	 branch_block_stmt_557/if_stmt_1035_dead_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_557/if_stmt_1035_eval_test/$entry
      -- CP-element group 116: 	 branch_block_stmt_557/if_stmt_1035_eval_test/$exit
      -- CP-element group 116: 	 branch_block_stmt_557/if_stmt_1035_eval_test/branch_req
      -- CP-element group 116: 	 branch_block_stmt_557/R_exitcond1_1036_place
      -- CP-element group 116: 	 branch_block_stmt_557/if_stmt_1035_if_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_557/if_stmt_1035_else_link/$entry
      -- 
    branch_req_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(116), ack => if_stmt_1035_branch_req_0); -- 
    sendB_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(115) & sendB_CP_1767_elements(103) & sendB_CP_1767_elements(99);
      gj_sendB_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  merge  transition  place  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	137 
    -- CP-element group 117:  members (13) 
      -- CP-element group 117: 	 branch_block_stmt_557/merge_stmt_1041__exit__
      -- CP-element group 117: 	 branch_block_stmt_557/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit
      -- CP-element group 117: 	 branch_block_stmt_557/if_stmt_1035_if_link/$exit
      -- CP-element group 117: 	 branch_block_stmt_557/if_stmt_1035_if_link/if_choice_transition
      -- CP-element group 117: 	 branch_block_stmt_557/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit
      -- CP-element group 117: 	 branch_block_stmt_557/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_557/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$exit
      -- CP-element group 117: 	 branch_block_stmt_557/merge_stmt_1041_PhiReqMerge
      -- CP-element group 117: 	 branch_block_stmt_557/merge_stmt_1041_PhiAck/$entry
      -- CP-element group 117: 	 branch_block_stmt_557/merge_stmt_1041_PhiAck/$exit
      -- CP-element group 117: 	 branch_block_stmt_557/merge_stmt_1041_PhiAck/dummy
      -- CP-element group 117: 	 branch_block_stmt_557/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_557/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1035_branch_ack_1, ack => sendB_CP_1767_elements(117)); -- 
    -- CP-element group 118:  fork  transition  place  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	132 
    -- CP-element group 118: 	133 
    -- CP-element group 118:  members (12) 
      -- CP-element group 118: 	 branch_block_stmt_557/if_stmt_1035_else_link/$exit
      -- CP-element group 118: 	 branch_block_stmt_557/if_stmt_1035_else_link/else_choice_transition
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/$entry
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/$entry
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/$entry
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/$entry
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1035_branch_ack_0, ack => sendB_CP_1767_elements(118)); -- 
    rr_3142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(118), ack => type_cast_984_inst_req_0); -- 
    cr_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(118), ack => type_cast_984_inst_req_1); -- 
    -- CP-element group 119:  transition  output  delay-element  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	1 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/phi_stmt_604/$exit
      -- CP-element group 119: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_608_konst_delay_trans
      -- CP-element group 119: 	 branch_block_stmt_557/bbx_xnph_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_req
      -- 
    phi_stmt_604_req_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_604_req_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(119), ack => phi_stmt_604_req_0); -- 
    -- Element group sendB_CP_1767_elements(119) is a control-delay.
    cp_element_119_delay: control_delay_element  generic map(name => " 119_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(1), ack => sendB_CP_1767_elements(119), clk => clk, reset =>reset);
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	50 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Sample/ra
      -- 
    ra_3023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_0, ack => sendB_CP_1767_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	50 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/Update/ca
      -- 
    ca_3028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_1, ack => sendB_CP_1767_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (6) 
      -- CP-element group 122: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/$exit
      -- CP-element group 122: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/$exit
      -- CP-element group 122: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_sources/type_cast_610/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_557/forx_xbody_forx_xbody_PhiReq/phi_stmt_604/phi_stmt_604_req
      -- 
    phi_stmt_604_req_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_604_req_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(122), ack => phi_stmt_604_req_1); -- 
    sendB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(120) & sendB_CP_1767_elements(121);
      gj_sendB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_557/merge_stmt_603_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_557/merge_stmt_603_PhiAck/$entry
      -- 
    sendB_CP_1767_elements(123) <= OrReduce(sendB_CP_1767_elements(119) & sendB_CP_1767_elements(122));
    -- CP-element group 124:  fork  transition  place  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	24 
    -- CP-element group 124: 	22 
    -- CP-element group 124: 	3 
    -- CP-element group 124: 	4 
    -- CP-element group 124: 	6 
    -- CP-element group 124: 	8 
    -- CP-element group 124: 	10 
    -- CP-element group 124: 	12 
    -- CP-element group 124: 	14 
    -- CP-element group 124: 	16 
    -- CP-element group 124: 	18 
    -- CP-element group 124: 	20 
    -- CP-element group 124:  members (53) 
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731__entry__
      -- CP-element group 124: 	 branch_block_stmt_557/merge_stmt_603__exit__
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/word_access_complete/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_update_start
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_resized_1
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_complete/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_scaled_1
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_665_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_scale_1/scale_rename_ack
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_scale_1/scale_rename_req
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Sample/req
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_scale_1/$exit
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Update/req
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_scale_1/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_resize_1/index_resize_ack
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_645_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_675_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_final_index_sum_regn_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_resize_1/index_resize_req
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_resize_1/$exit
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_resize_1/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/array_obj_ref_616_index_computed_1
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_655_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/word_access_complete/word_0/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/ptr_deref_621_Update/word_access_complete/word_0/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/addr_of_617_complete/req
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_635_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_625_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_685_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_update_start_
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_557/assign_stmt_618_to_assign_stmt_731/type_cast_695_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_557/merge_stmt_603_PhiAck/$exit
      -- CP-element group 124: 	 branch_block_stmt_557/merge_stmt_603_PhiAck/phi_stmt_604_ack
      -- 
    phi_stmt_604_ack_3034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_604_ack_0, ack => sendB_CP_1767_elements(124)); -- 
    cr_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_625_inst_req_1); -- 
    cr_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_675_inst_req_1); -- 
    cr_2013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_665_inst_req_1); -- 
    cr_1971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_635_inst_req_1); -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => array_obj_ref_616_index_offset_req_0); -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => array_obj_ref_616_index_offset_req_1); -- 
    cr_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_645_inst_req_1); -- 
    cr_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_655_inst_req_1); -- 
    cr_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => ptr_deref_621_load_0_req_1); -- 
    req_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => addr_of_617_final_reg_req_1); -- 
    cr_2041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_685_inst_req_1); -- 
    cr_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(124), ack => type_cast_695_inst_req_1); -- 
    -- CP-element group 125:  transition  output  delay-element  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	2 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/$exit
      -- CP-element group 125: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/phi_stmt_764/$exit
      -- CP-element group 125: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_768_konst_delay_trans
      -- CP-element group 125: 	 branch_block_stmt_557/entry_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_req
      -- 
    phi_stmt_764_req_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_764_req_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(125), ack => phi_stmt_764_req_0); -- 
    -- Element group sendB_CP_1767_elements(125) is a control-delay.
    cp_element_125_delay: control_delay_element  generic map(name => " 125_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(2), ack => sendB_CP_1767_elements(125), clk => clk, reset =>reset);
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	49 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Sample/ra
      -- 
    ra_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_770_inst_ack_0, ack => sendB_CP_1767_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	49 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/Update/ca
      -- 
    ca_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_770_inst_ack_1, ack => sendB_CP_1767_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 128: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/$exit
      -- CP-element group 128: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/$exit
      -- CP-element group 128: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_557/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_764/phi_stmt_764_req
      -- 
    phi_stmt_764_req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_764_req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(128), ack => phi_stmt_764_req_1); -- 
    sendB_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(127) & sendB_CP_1767_elements(126);
      gj_sendB_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  merge  transition  place  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: 	125 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_557/merge_stmt_763_PhiReqMerge
      -- CP-element group 129: 	 branch_block_stmt_557/merge_stmt_763_PhiAck/$entry
      -- 
    sendB_CP_1767_elements(129) <= OrReduce(sendB_CP_1767_elements(128) & sendB_CP_1767_elements(125));
    -- CP-element group 130:  branch  transition  place  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	51 
    -- CP-element group 130: 	52 
    -- CP-element group 130:  members (15) 
      -- CP-element group 130: 	 branch_block_stmt_557/merge_stmt_763__exit__
      -- CP-element group 130: 	 branch_block_stmt_557/if_stmt_784__entry__
      -- CP-element group 130: 	 branch_block_stmt_557/assign_stmt_777_to_assign_stmt_783__exit__
      -- CP-element group 130: 	 branch_block_stmt_557/assign_stmt_777_to_assign_stmt_783__entry__
      -- CP-element group 130: 	 branch_block_stmt_557/assign_stmt_777_to_assign_stmt_783/$entry
      -- CP-element group 130: 	 branch_block_stmt_557/assign_stmt_777_to_assign_stmt_783/$exit
      -- CP-element group 130: 	 branch_block_stmt_557/if_stmt_784_dead_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_557/if_stmt_784_eval_test/$entry
      -- CP-element group 130: 	 branch_block_stmt_557/if_stmt_784_eval_test/$exit
      -- CP-element group 130: 	 branch_block_stmt_557/if_stmt_784_eval_test/branch_req
      -- CP-element group 130: 	 branch_block_stmt_557/R_tobool_785_place
      -- CP-element group 130: 	 branch_block_stmt_557/if_stmt_784_if_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_557/if_stmt_784_else_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_557/merge_stmt_763_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_557/merge_stmt_763_PhiAck/phi_stmt_764_ack
      -- 
    phi_stmt_764_ack_3088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_764_ack_0, ack => sendB_CP_1767_elements(130)); -- 
    branch_req_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(130), ack => if_stmt_784_branch_req_0); -- 
    -- CP-element group 131:  transition  output  delay-element  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	98 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	135 
    -- CP-element group 131:  members (5) 
      -- CP-element group 131: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- CP-element group 131: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/$exit
      -- CP-element group 131: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/$exit
      -- CP-element group 131: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_982_konst_delay_trans
      -- CP-element group 131: 	 branch_block_stmt_557/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_req
      -- 
    phi_stmt_978_req_3123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_978_req_3123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(131), ack => phi_stmt_978_req_0); -- 
    -- Element group sendB_CP_1767_elements(131) is a control-delay.
    cp_element_131_delay: control_delay_element  generic map(name => " 131_delay", delay_value => 1)  port map(req => sendB_CP_1767_elements(98), ack => sendB_CP_1767_elements(131), clk => clk, reset =>reset);
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	118 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Sample/ra
      -- 
    ra_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_984_inst_ack_0, ack => sendB_CP_1767_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	118 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/Update/ca
      -- 
    ca_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_984_inst_ack_1, ack => sendB_CP_1767_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- CP-element group 134: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/$exit
      -- CP-element group 134: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/$exit
      -- CP-element group 134: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/$exit
      -- CP-element group 134: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_sources/type_cast_984/SplitProtocol/$exit
      -- CP-element group 134: 	 branch_block_stmt_557/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_978/phi_stmt_978_req
      -- 
    phi_stmt_978_req_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_978_req_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(134), ack => phi_stmt_978_req_1); -- 
    sendB_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1767_elements(132) & sendB_CP_1767_elements(133);
      gj_sendB_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1767_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  merge  transition  place  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	131 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_557/merge_stmt_977_PhiReqMerge
      -- CP-element group 135: 	 branch_block_stmt_557/merge_stmt_977_PhiAck/$entry
      -- 
    sendB_CP_1767_elements(135) <= OrReduce(sendB_CP_1767_elements(131) & sendB_CP_1767_elements(134));
    -- CP-element group 136:  fork  transition  place  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	108 
    -- CP-element group 136: 	102 
    -- CP-element group 136: 	100 
    -- CP-element group 136: 	106 
    -- CP-element group 136: 	103 
    -- CP-element group 136: 	104 
    -- CP-element group 136: 	112 
    -- CP-element group 136: 	99 
    -- CP-element group 136:  members (53) 
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Update/req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Update/req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/merge_stmt_977__exit__
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034__entry__
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_update_start_
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_final_index_sum_regn_update_start
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_complete/req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_final_index_sum_regn_update_start
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_scale_1/scale_rename_ack
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_scale_1/scale_rename_req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_scale_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_scale_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_resize_1/index_resize_ack
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_resize_1/index_resize_req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_resize_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_resize_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_computed_1
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_scaled_1
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_scale_1/scale_rename_ack
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_scale_1/scale_rename_req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_index_resized_1
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_scale_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_scale_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_update_start_
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_update_start_
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_resize_1/index_resize_ack
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_resize_1/index_resize_req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_resize_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_complete/req
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_resize_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_computed_1
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/word_access_complete/word_0/cr
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_scaled_1
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/word_access_complete/word_0/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_1008_index_resized_1
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1012_Update/word_access_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/array_obj_ref_996_update_start_
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/word_access_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/word_access_complete/word_0/$entry
      -- CP-element group 136: 	 branch_block_stmt_557/assign_stmt_991_to_assign_stmt_1034/ptr_deref_1019_Update/word_access_complete/word_0/cr
      -- CP-element group 136: 	 branch_block_stmt_557/merge_stmt_977_PhiAck/$exit
      -- CP-element group 136: 	 branch_block_stmt_557/merge_stmt_977_PhiAck/phi_stmt_978_ack
      -- 
    phi_stmt_978_ack_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_978_ack_0, ack => sendB_CP_1767_elements(136)); -- 
    req_2817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => array_obj_ref_1008_index_offset_req_1); -- 
    req_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => array_obj_ref_996_index_offset_req_1); -- 
    req_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => array_obj_ref_1008_index_offset_req_0); -- 
    req_2785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => array_obj_ref_996_final_reg_req_1); -- 
    req_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => array_obj_ref_996_index_offset_req_0); -- 
    req_2832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => array_obj_ref_1008_final_reg_req_1); -- 
    cr_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => ptr_deref_1012_load_0_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1767_elements(136), ack => ptr_deref_1019_load_0_req_1); -- 
    -- CP-element group 137:  merge  transition  place  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	117 
    -- CP-element group 137: 	97 
    -- CP-element group 137: 	51 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (16) 
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1043__exit__
      -- CP-element group 137: 	 branch_block_stmt_557/branch_block_stmt_557__exit__
      -- CP-element group 137: 	 branch_block_stmt_557/$exit
      -- CP-element group 137: 	 $exit
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1045__exit__
      -- CP-element group 137: 	 branch_block_stmt_557/return__
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1045_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1043_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1043_PhiAck/$entry
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1043_PhiAck/$exit
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1043_PhiAck/dummy
      -- CP-element group 137: 	 branch_block_stmt_557/return___PhiReq/$entry
      -- CP-element group 137: 	 branch_block_stmt_557/return___PhiReq/$exit
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1045_PhiAck/$entry
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1045_PhiAck/$exit
      -- CP-element group 137: 	 branch_block_stmt_557/merge_stmt_1045_PhiAck/dummy
      -- 
    sendB_CP_1767_elements(137) <= OrReduce(sendB_CP_1767_elements(117) & sendB_CP_1767_elements(97) & sendB_CP_1767_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_759_wire : std_logic_vector(63 downto 0);
    signal R_indvar_615_resized : std_logic_vector(13 downto 0);
    signal R_indvar_615_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_798_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_798_scaled : std_logic_vector(13 downto 0);
    signal R_tmp2_995_resized : std_logic_vector(2 downto 0);
    signal R_tmp2_995_scaled : std_logic_vector(2 downto 0);
    signal R_tmp3_1007_resized : std_logic_vector(2 downto 0);
    signal R_tmp3_1007_scaled : std_logic_vector(2 downto 0);
    signal and70_777 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1008_constant_part_of_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1008_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1008_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1008_offset_scale_factor_1 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1008_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1008_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_616_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_616_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_616_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_616_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_616_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_616_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_799_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_799_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_799_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_799_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_799_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_799_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_996_constant_part_of_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_996_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_996_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_996_offset_scale_factor_1 : std_logic_vector(2 downto 0);
    signal array_obj_ref_996_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_996_root_address : std_logic_vector(2 downto 0);
    signal arrayidx11x_xi_843 : std_logic_vector(31 downto 0);
    signal arrayidx17x_xi_864 : std_logic_vector(31 downto 0);
    signal arrayidx23x_xi_885 : std_logic_vector(31 downto 0);
    signal arrayidx29x_xi_906 : std_logic_vector(31 downto 0);
    signal arrayidx35x_xi_927 : std_logic_vector(31 downto 0);
    signal arrayidx43x_xi_997 : std_logic_vector(31 downto 0);
    signal arrayidx48x_xi_1009 : std_logic_vector(31 downto 0);
    signal arrayidx5x_xi_822 : std_logic_vector(31 downto 0);
    signal arrayidx_618 : std_logic_vector(31 downto 0);
    signal arrayidxx_xi_801 : std_logic_vector(31 downto 0);
    signal cmp53x_xi_937 : std_logic_vector(0 downto 0);
    signal cmp77_569 : std_logic_vector(0 downto 0);
    signal conv10x_xi_836 : std_logic_vector(7 downto 0);
    signal conv14_636 : std_logic_vector(7 downto 0);
    signal conv16x_xi_857 : std_logic_vector(7 downto 0);
    signal conv20_646 : std_logic_vector(7 downto 0);
    signal conv22x_xi_878 : std_logic_vector(7 downto 0);
    signal conv26_656 : std_logic_vector(7 downto 0);
    signal conv28x_xi_899 : std_logic_vector(7 downto 0);
    signal conv32_666 : std_logic_vector(7 downto 0);
    signal conv34x_xi_920 : std_logic_vector(7 downto 0);
    signal conv38_676 : std_logic_vector(7 downto 0);
    signal conv44_686 : std_logic_vector(7 downto 0);
    signal conv50_696 : std_logic_vector(7 downto 0);
    signal conv74_794 : std_logic_vector(15 downto 0);
    signal conv8_626 : std_logic_vector(7 downto 0);
    signal convx_xi_815 : std_logic_vector(7 downto 0);
    signal exitcond1_1034 : std_logic_vector(0 downto 0);
    signal exitcond_731 : std_logic_vector(0 downto 0);
    signal iNsTr_29_962 : std_logic_vector(63 downto 0);
    signal indvar_604 : std_logic_vector(63 downto 0);
    signal indvarx_xi_978 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_726 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi_1029 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_764 : std_logic_vector(63 downto 0);
    signal out_datax_xi_563 : std_logic_vector(31 downto 0);
    signal phitmp_761 : std_logic_vector(63 downto 0);
    signal ptr_deref_1012_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1012_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1012_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1012_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1012_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1019_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1019_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1019_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1019_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1019_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_621_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_621_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_621_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_621_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_621_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_804_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_804_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_804_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_804_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_804_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_824_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_824_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_824_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_824_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_824_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_824_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_845_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_845_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_845_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_845_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_845_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_845_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_866_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_866_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_866_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_866_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_866_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_866_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_887_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_887_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_887_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_887_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_887_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_887_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_908_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_908_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_908_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_908_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_908_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_908_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_929_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_929_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_929_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_929_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_929_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_929_word_offset_0 : std_logic_vector(2 downto 0);
    signal shr11_632 : std_logic_vector(63 downto 0);
    signal shr13x_xi_853 : std_logic_vector(63 downto 0);
    signal shr17_642 : std_logic_vector(63 downto 0);
    signal shr19x_xi_874 : std_logic_vector(63 downto 0);
    signal shr23_652 : std_logic_vector(63 downto 0);
    signal shr25x_xi_895 : std_logic_vector(63 downto 0);
    signal shr29_662 : std_logic_vector(63 downto 0);
    signal shr31x_xi_916 : std_logic_vector(63 downto 0);
    signal shr35_672 : std_logic_vector(63 downto 0);
    signal shr41_682 : std_logic_vector(63 downto 0);
    signal shr47_692 : std_logic_vector(63 downto 0);
    signal shr7x_xi_832 : std_logic_vector(63 downto 0);
    signal shr_582 : std_logic_vector(63 downto 0);
    signal shrx_xi_811 : std_logic_vector(63 downto 0);
    signal tmp1x_xi_805 : std_logic_vector(63 downto 0);
    signal tmp2_991 : std_logic_vector(63 downto 0);
    signal tmp3_1003 : std_logic_vector(63 downto 0);
    signal tmp44x_xi_1013 : std_logic_vector(7 downto 0);
    signal tmp49x_xi_1020 : std_logic_vector(7 downto 0);
    signal tmp55x_xi_950 : std_logic_vector(0 downto 0);
    signal tmp58x_xi_975 : std_logic_vector(63 downto 0);
    signal tmp5_622 : std_logic_vector(63 downto 0);
    signal tmp80_588 : std_logic_vector(0 downto 0);
    signal tmp81_751 : std_logic_vector(63 downto 0);
    signal tmp_594 : std_logic_vector(0 downto 0);
    signal tmpx_xopx_xi_956 : std_logic_vector(63 downto 0);
    signal tobool_783 : std_logic_vector(0 downto 0);
    signal type_cast_1001_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1027_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_580_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_586_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_592_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_599_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_608_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_610_wire : std_logic_vector(63 downto 0);
    signal type_cast_630_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_640_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_650_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_660_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_670_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_680_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_690_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_743_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_749_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire : std_logic_vector(63 downto 0);
    signal type_cast_758_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_768_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_770_wire : std_logic_vector(63 downto 0);
    signal type_cast_775_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_781_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_830_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_851_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_872_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_914_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_935_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_954_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_960_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_966_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_973_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_982_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_984_wire : std_logic_vector(63 downto 0);
    signal type_cast_989_wire_constant : std_logic_vector(63 downto 0);
    signal umax4_601 : std_logic_vector(63 downto 0);
    signal umax_745 : std_logic_vector(63 downto 0);
    signal xx_xopx_xi_968 : std_logic_vector(63 downto 0);
    signal xxsendBxxbodyxxout_datax_xi_alloc_base_address : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    array_obj_ref_1008_constant_part_of_offset <= "000";
    array_obj_ref_1008_offset_scale_factor_0 <= "110";
    array_obj_ref_1008_offset_scale_factor_1 <= "001";
    array_obj_ref_1008_resized_base_address <= "000";
    array_obj_ref_616_constant_part_of_offset <= "00000000000000";
    array_obj_ref_616_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_616_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_616_resized_base_address <= "00000000000000";
    array_obj_ref_799_constant_part_of_offset <= "00000000000000";
    array_obj_ref_799_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_799_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_799_resized_base_address <= "00000000000000";
    array_obj_ref_996_constant_part_of_offset <= "000";
    array_obj_ref_996_offset_scale_factor_0 <= "110";
    array_obj_ref_996_offset_scale_factor_1 <= "001";
    array_obj_ref_996_resized_base_address <= "000";
    arrayidx11x_xi_843 <= "00000000000000000000000000000100";
    arrayidx17x_xi_864 <= "00000000000000000000000000000011";
    arrayidx23x_xi_885 <= "00000000000000000000000000000010";
    arrayidx29x_xi_906 <= "00000000000000000000000000000001";
    arrayidx35x_xi_927 <= "00000000000000000000000000000000";
    arrayidx5x_xi_822 <= "00000000000000000000000000000101";
    out_datax_xi_563 <= "00000000000000000000000000000000";
    ptr_deref_1012_word_offset_0 <= "000";
    ptr_deref_1019_word_offset_0 <= "000";
    ptr_deref_621_word_offset_0 <= "00000000000000";
    ptr_deref_804_word_offset_0 <= "00000000000000";
    ptr_deref_824_word_offset_0 <= "000";
    ptr_deref_845_word_offset_0 <= "000";
    ptr_deref_866_word_offset_0 <= "000";
    ptr_deref_887_word_offset_0 <= "000";
    ptr_deref_908_word_offset_0 <= "000";
    ptr_deref_929_word_offset_0 <= "000";
    type_cast_1001_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1027_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_567_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_580_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_586_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_592_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_599_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_608_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_630_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_640_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_650_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_660_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_670_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_680_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_690_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_743_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_749_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_758_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_768_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_775_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_781_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_809_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_830_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_851_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_872_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_893_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_914_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_935_wire_constant <= "0000000000000000";
    type_cast_948_wire_constant <= "0000000000000001";
    type_cast_954_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_960_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_966_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_973_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_982_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_989_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    xxsendBxxbodyxxout_datax_xi_alloc_base_address <= "000";
    phi_stmt_604: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_608_wire_constant & type_cast_610_wire;
      req <= phi_stmt_604_req_0 & phi_stmt_604_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_604",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_604_ack_0,
          idata => idata,
          odata => indvar_604,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_604
    phi_stmt_764: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_768_wire_constant & type_cast_770_wire;
      req <= phi_stmt_764_req_0 & phi_stmt_764_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_764",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_764_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_764,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_764
    phi_stmt_978: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_982_wire_constant & type_cast_984_wire;
      req <= phi_stmt_978_req_0 & phi_stmt_978_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_978",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_978_ack_0,
          idata => idata,
          odata => indvarx_xi_978,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_978
    -- flow-through select operator MUX_600_inst
    umax4_601 <= shr_582 when (tmp_594(0) /=  '0') else type_cast_599_wire_constant;
    -- flow-through select operator MUX_744_inst
    umax_745 <= shr_582 when (tmp80_588(0) /=  '0') else type_cast_743_wire_constant;
    -- flow-through select operator MUX_974_inst
    tmp58x_xi_975 <= xx_xopx_xi_968 when (tmp55x_xi_950(0) /=  '0') else type_cast_973_wire_constant;
    addr_of_617_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_617_final_reg_req_0;
      addr_of_617_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_617_final_reg_req_1;
      addr_of_617_final_reg_ack_1<= rack(0);
      addr_of_617_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_617_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_616_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_800_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_800_final_reg_req_0;
      addr_of_800_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_800_final_reg_req_1;
      addr_of_800_final_reg_ack_1<= rack(0);
      addr_of_800_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_800_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_799_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidxx_xi_801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    array_obj_ref_1008_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= array_obj_ref_1008_final_reg_req_0;
      array_obj_ref_1008_final_reg_ack_0<= wack(0);
      rreq(0) <= array_obj_ref_1008_final_reg_req_1;
      array_obj_ref_1008_final_reg_ack_1<= rack(0);
      array_obj_ref_1008_final_reg : InterlockBuffer generic map ( -- 
        name => "array_obj_ref_1008_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1008_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx48x_xi_1009,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    array_obj_ref_996_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= array_obj_ref_996_final_reg_req_0;
      array_obj_ref_996_final_reg_ack_0<= wack(0);
      rreq(0) <= array_obj_ref_996_final_reg_req_1;
      array_obj_ref_996_final_reg_ack_1<= rack(0);
      array_obj_ref_996_final_reg : InterlockBuffer generic map ( -- 
        name => "array_obj_ref_996_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_996_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx43x_xi_997,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_610_inst_req_0;
      type_cast_610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_610_inst_req_1;
      type_cast_610_inst_ack_1<= rack(0);
      type_cast_610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_610_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_625_inst_req_0;
      type_cast_625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_625_inst_req_1;
      type_cast_625_inst_ack_1<= rack(0);
      type_cast_625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_626,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_635_inst_req_0;
      type_cast_635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_635_inst_req_1;
      type_cast_635_inst_ack_1<= rack(0);
      type_cast_635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr11_632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_645_inst_req_0;
      type_cast_645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_645_inst_req_1;
      type_cast_645_inst_ack_1<= rack(0);
      type_cast_645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_645_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_655_inst_req_0;
      type_cast_655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_655_inst_req_1;
      type_cast_655_inst_ack_1<= rack(0);
      type_cast_655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_652,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_665_inst_req_0;
      type_cast_665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_665_inst_req_1;
      type_cast_665_inst_ack_1<= rack(0);
      type_cast_665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_662,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_675_inst_req_0;
      type_cast_675_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_675_inst_req_1;
      type_cast_675_inst_ack_1<= rack(0);
      type_cast_675_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_675_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_676,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_685_inst_req_0;
      type_cast_685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_685_inst_req_1;
      type_cast_685_inst_ack_1<= rack(0);
      type_cast_685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_682,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_695_inst_req_0;
      type_cast_695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_695_inst_req_1;
      type_cast_695_inst_ack_1<= rack(0);
      type_cast_695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_755_inst
    process(tmp81_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp81_751(63 downto 0);
      type_cast_755_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_760_inst
    process(ASHR_i64_i64_759_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_759_wire(63 downto 0);
      phitmp_761 <= tmp_var; -- 
    end process;
    type_cast_770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_770_inst_req_0;
      type_cast_770_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_770_inst_req_1;
      type_cast_770_inst_ack_1<= rack(0);
      type_cast_770_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_770_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_793_inst_req_0;
      type_cast_793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_793_inst_req_1;
      type_cast_793_inst_ack_1<= rack(0);
      type_cast_793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => and70_777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_814_inst_req_0;
      type_cast_814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_814_inst_req_1;
      type_cast_814_inst_ack_1<= rack(0);
      type_cast_814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_814_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xi_811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_835_inst_req_0;
      type_cast_835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_835_inst_req_1;
      type_cast_835_inst_ack_1<= rack(0);
      type_cast_835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr7x_xi_832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10x_xi_836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_856_inst_req_0;
      type_cast_856_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_856_inst_req_1;
      type_cast_856_inst_ack_1<= rack(0);
      type_cast_856_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_856_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr13x_xi_853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16x_xi_857,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_877_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_877_inst_req_0;
      type_cast_877_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_877_inst_req_1;
      type_cast_877_inst_ack_1<= rack(0);
      type_cast_877_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_877_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr19x_xi_874,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22x_xi_878,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_898_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_898_inst_req_0;
      type_cast_898_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_898_inst_req_1;
      type_cast_898_inst_ack_1<= rack(0);
      type_cast_898_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_898_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr25x_xi_895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28x_xi_899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_919_inst_req_0;
      type_cast_919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_919_inst_req_1;
      type_cast_919_inst_ack_1<= rack(0);
      type_cast_919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr31x_xi_916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34x_xi_920,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_984_inst_req_0;
      type_cast_984_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_984_inst_req_1;
      type_cast_984_inst_ack_1<= rack(0);
      type_cast_984_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_984_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1008_index_1_rename
    process(R_tmp3_1007_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp3_1007_resized;
      ov(2 downto 0) := iv;
      R_tmp3_1007_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1008_index_1_resize
    process(tmp3_1003) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp3_1003;
      ov := iv(2 downto 0);
      R_tmp3_1007_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1008_root_address_inst
    process(array_obj_ref_1008_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1008_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_1008_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_616_index_1_rename
    process(R_indvar_615_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_615_resized;
      ov(13 downto 0) := iv;
      R_indvar_615_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_616_index_1_resize
    process(indvar_604) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_604;
      ov := iv(13 downto 0);
      R_indvar_615_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_616_root_address_inst
    process(array_obj_ref_616_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_616_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_616_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_799_index_1_rename
    process(R_ix_x0x_xlcssa_798_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_798_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_798_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_799_index_1_resize
    process(ix_x0x_xlcssa_764) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_764;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_798_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_799_root_address_inst
    process(array_obj_ref_799_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_799_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_799_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_996_index_1_rename
    process(R_tmp2_995_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp2_995_resized;
      ov(2 downto 0) := iv;
      R_tmp2_995_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_996_index_1_resize
    process(tmp2_991) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp2_991;
      ov := iv(2 downto 0);
      R_tmp2_995_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_996_root_address_inst
    process(array_obj_ref_996_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_996_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_996_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1012_addr_0
    process(ptr_deref_1012_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1012_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1012_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1012_base_resize
    process(arrayidx43x_xi_997) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx43x_xi_997;
      ov := iv(2 downto 0);
      ptr_deref_1012_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1012_gather_scatter
    process(ptr_deref_1012_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1012_data_0;
      ov(7 downto 0) := iv;
      tmp44x_xi_1013 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1012_root_address_inst
    process(ptr_deref_1012_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1012_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1012_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_addr_0
    process(ptr_deref_1019_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1019_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1019_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_base_resize
    process(arrayidx48x_xi_1009) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx48x_xi_1009;
      ov := iv(2 downto 0);
      ptr_deref_1019_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_gather_scatter
    process(ptr_deref_1019_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1019_data_0;
      ov(7 downto 0) := iv;
      tmp49x_xi_1020 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_root_address_inst
    process(ptr_deref_1019_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1019_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1019_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_621_addr_0
    process(ptr_deref_621_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_621_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_621_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_621_base_resize
    process(arrayidx_618) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_618;
      ov := iv(13 downto 0);
      ptr_deref_621_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_621_gather_scatter
    process(ptr_deref_621_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_621_data_0;
      ov(63 downto 0) := iv;
      tmp5_622 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_621_root_address_inst
    process(ptr_deref_621_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_621_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_621_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_addr_0
    process(ptr_deref_804_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_804_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_804_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_base_resize
    process(arrayidxx_xi_801) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidxx_xi_801;
      ov := iv(13 downto 0);
      ptr_deref_804_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_gather_scatter
    process(ptr_deref_804_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_804_data_0;
      ov(63 downto 0) := iv;
      tmp1x_xi_805 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_root_address_inst
    process(ptr_deref_804_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_804_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_804_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_addr_0
    process(ptr_deref_824_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_824_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_824_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_base_resize
    process(arrayidx5x_xi_822) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx5x_xi_822;
      ov := iv(2 downto 0);
      ptr_deref_824_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_gather_scatter
    process(convx_xi_815) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := convx_xi_815;
      ov(7 downto 0) := iv;
      ptr_deref_824_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_root_address_inst
    process(ptr_deref_824_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_824_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_824_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_845_addr_0
    process(ptr_deref_845_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_845_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_845_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_845_base_resize
    process(arrayidx11x_xi_843) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx11x_xi_843;
      ov := iv(2 downto 0);
      ptr_deref_845_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_845_gather_scatter
    process(conv10x_xi_836) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv10x_xi_836;
      ov(7 downto 0) := iv;
      ptr_deref_845_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_845_root_address_inst
    process(ptr_deref_845_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_845_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_845_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_866_addr_0
    process(ptr_deref_866_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_866_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_866_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_866_base_resize
    process(arrayidx17x_xi_864) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx17x_xi_864;
      ov := iv(2 downto 0);
      ptr_deref_866_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_866_gather_scatter
    process(conv16x_xi_857) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16x_xi_857;
      ov(7 downto 0) := iv;
      ptr_deref_866_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_866_root_address_inst
    process(ptr_deref_866_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_866_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_866_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_887_addr_0
    process(ptr_deref_887_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_887_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_887_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_887_base_resize
    process(arrayidx23x_xi_885) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx23x_xi_885;
      ov := iv(2 downto 0);
      ptr_deref_887_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_887_gather_scatter
    process(conv22x_xi_878) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv22x_xi_878;
      ov(7 downto 0) := iv;
      ptr_deref_887_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_887_root_address_inst
    process(ptr_deref_887_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_887_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_887_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_908_addr_0
    process(ptr_deref_908_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_908_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_908_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_908_base_resize
    process(arrayidx29x_xi_906) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx29x_xi_906;
      ov := iv(2 downto 0);
      ptr_deref_908_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_908_gather_scatter
    process(conv28x_xi_899) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv28x_xi_899;
      ov(7 downto 0) := iv;
      ptr_deref_908_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_908_root_address_inst
    process(ptr_deref_908_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_908_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_908_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_addr_0
    process(ptr_deref_929_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_929_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_929_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_base_resize
    process(arrayidx35x_xi_927) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx35x_xi_927;
      ov := iv(2 downto 0);
      ptr_deref_929_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_gather_scatter
    process(conv34x_xi_920) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv34x_xi_920;
      ov(7 downto 0) := iv;
      ptr_deref_929_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_root_address_inst
    process(ptr_deref_929_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_929_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_929_root_address <= ov(2 downto 0);
      --
    end process;
    if_stmt_1035_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1034;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1035_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1035_branch_req_0,
          ack0 => if_stmt_1035_branch_ack_0,
          ack1 => if_stmt_1035_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_570_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_569;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_570_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_570_branch_req_0,
          ack0 => if_stmt_570_branch_ack_0,
          ack1 => if_stmt_570_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_732_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_731;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_732_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_732_branch_req_0,
          ack0 => if_stmt_732_branch_ack_0,
          ack1 => if_stmt_732_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_784_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_783;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_784_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_784_branch_req_0,
          ack0 => if_stmt_784_branch_ack_0,
          ack1 => if_stmt_784_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_938_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp53x_xi_937;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_938_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_938_branch_req_0,
          ack0 => if_stmt_938_branch_ack_0,
          ack1 => if_stmt_938_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1002_inst
    process(tmp2_991) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_991, type_cast_1001_wire_constant, tmp_var);
      tmp3_1003 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1028_inst
    process(indvarx_xi_978) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvarx_xi_978, type_cast_1027_wire_constant, tmp_var);
      indvarx_xnextx_xi_1029 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_725_inst
    process(indvar_604) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_604, type_cast_724_wire_constant, tmp_var);
      indvarx_xnext_726 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_955_inst
    process(and70_777) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(and70_777, type_cast_954_wire_constant, tmp_var);
      tmpx_xopx_xi_956 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_967_inst
    process(iNsTr_29_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_29_962, type_cast_966_wire_constant, tmp_var);
      xx_xopx_xi_968 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_776_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(size_buffer, type_cast_775_wire_constant, tmp_var);
      and70_777 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_961_inst
    process(tmpx_xopx_xi_956) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tmpx_xopx_xi_956, type_cast_960_wire_constant, tmp_var);
      iNsTr_29_962 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_759_inst
    process(type_cast_755_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_755_wire, type_cast_758_wire_constant, tmp_var);
      ASHR_i64_i64_759_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_936_inst
    process(conv74_794) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_794, type_cast_935_wire_constant, tmp_var);
      cmp53x_xi_937 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1033_inst
    process(indvarx_xnextx_xi_1029, tmp58x_xi_975) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnextx_xi_1029, tmp58x_xi_975, tmp_var);
      exitcond1_1034 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_730_inst
    process(indvarx_xnext_726, umax4_601) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_726, umax4_601, tmp_var);
      exitcond_731 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_782_inst
    process(and70_777) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and70_777, type_cast_781_wire_constant, tmp_var);
      tobool_783 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_581_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_580_wire_constant, tmp_var);
      shr_582 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_631_inst
    process(tmp5_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_622, type_cast_630_wire_constant, tmp_var);
      shr11_632 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_641_inst
    process(tmp5_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_622, type_cast_640_wire_constant, tmp_var);
      shr17_642 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_651_inst
    process(tmp5_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_622, type_cast_650_wire_constant, tmp_var);
      shr23_652 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_661_inst
    process(tmp5_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_622, type_cast_660_wire_constant, tmp_var);
      shr29_662 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_671_inst
    process(tmp5_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_622, type_cast_670_wire_constant, tmp_var);
      shr35_672 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_681_inst
    process(tmp5_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_622, type_cast_680_wire_constant, tmp_var);
      shr41_682 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_691_inst
    process(tmp5_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_622, type_cast_690_wire_constant, tmp_var);
      shr47_692 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_810_inst
    process(tmp1x_xi_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_805, type_cast_809_wire_constant, tmp_var);
      shrx_xi_811 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_831_inst
    process(tmp1x_xi_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_805, type_cast_830_wire_constant, tmp_var);
      shr7x_xi_832 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_852_inst
    process(tmp1x_xi_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_805, type_cast_851_wire_constant, tmp_var);
      shr13x_xi_853 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_873_inst
    process(tmp1x_xi_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_805, type_cast_872_wire_constant, tmp_var);
      shr19x_xi_874 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_894_inst
    process(tmp1x_xi_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_805, type_cast_893_wire_constant, tmp_var);
      shr25x_xi_895 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_915_inst
    process(tmp1x_xi_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_805, type_cast_914_wire_constant, tmp_var);
      shr31x_xi_916 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_990_inst
    process(indvarx_xi_978) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvarx_xi_978, type_cast_989_wire_constant, tmp_var);
      tmp2_991 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_750_inst
    process(umax_745) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_745, type_cast_749_wire_constant, tmp_var);
      tmp81_751 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_949_inst
    process(conv74_794) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv74_794, type_cast_948_wire_constant, tmp_var);
      tmp55x_xi_950 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_568_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_567_wire_constant, tmp_var);
      cmp77_569 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_587_inst
    process(shr_582) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_582, type_cast_586_wire_constant, tmp_var);
      tmp80_588 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_593_inst
    process(shr_582) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_582, type_cast_592_wire_constant, tmp_var);
      tmp_594 <= tmp_var; --
    end process;
    -- shared split operator group (32) : array_obj_ref_1008_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_tmp3_1007_scaled;
      array_obj_ref_1008_final_offset <= data_out(2 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1008_index_offset_req_0;
      array_obj_ref_1008_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1008_index_offset_req_1;
      array_obj_ref_1008_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : array_obj_ref_616_index_offset 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_615_scaled;
      array_obj_ref_616_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_616_index_offset_req_0;
      array_obj_ref_616_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_616_index_offset_req_1;
      array_obj_ref_616_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : array_obj_ref_799_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_798_scaled;
      array_obj_ref_799_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_799_index_offset_req_0;
      array_obj_ref_799_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_799_index_offset_req_1;
      array_obj_ref_799_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_996_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_tmp2_995_scaled;
      array_obj_ref_996_final_offset <= data_out(2 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_996_index_offset_req_0;
      array_obj_ref_996_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_996_index_offset_req_1;
      array_obj_ref_996_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared load operator group (0) : ptr_deref_1012_load_0 ptr_deref_1019_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1012_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1019_load_0_req_0;
      ptr_deref_1012_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1019_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1012_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1019_load_0_req_1;
      ptr_deref_1012_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1019_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1012_word_address_0 & ptr_deref_1019_word_address_0;
      ptr_deref_1012_data_0 <= data_out(15 downto 8);
      ptr_deref_1019_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 3,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(2 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_621_load_0 ptr_deref_804_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_621_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_804_load_0_req_0;
      ptr_deref_621_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_804_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_621_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_804_load_0_req_1;
      ptr_deref_621_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_804_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_621_word_address_0 & ptr_deref_804_word_address_0;
      ptr_deref_621_data_0 <= data_out(127 downto 64);
      ptr_deref_804_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_929_store_0 ptr_deref_824_store_0 ptr_deref_845_store_0 ptr_deref_866_store_0 ptr_deref_887_store_0 ptr_deref_908_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(17 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_929_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_824_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_845_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_866_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_887_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_908_store_0_req_0;
      ptr_deref_929_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_824_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_845_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_866_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_887_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_908_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_929_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_824_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_845_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_866_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_887_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_908_store_0_req_1;
      ptr_deref_929_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_824_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_845_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_866_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_887_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_908_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_929_word_address_0 & ptr_deref_824_word_address_0 & ptr_deref_845_word_address_0 & ptr_deref_866_word_address_0 & ptr_deref_887_word_address_0 & ptr_deref_908_word_address_0;
      data_in <= ptr_deref_929_data_0 & ptr_deref_824_data_0 & ptr_deref_845_data_0 & ptr_deref_866_data_0 & ptr_deref_887_data_0 & ptr_deref_908_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 3,
        data_width => 8,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(2 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 6,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1014_inst WPIPE_maxpool_output_pipe_697_inst WPIPE_maxpool_output_pipe_700_inst WPIPE_maxpool_output_pipe_703_inst WPIPE_maxpool_output_pipe_706_inst WPIPE_maxpool_output_pipe_709_inst WPIPE_maxpool_output_pipe_712_inst WPIPE_maxpool_output_pipe_715_inst WPIPE_maxpool_output_pipe_718_inst WPIPE_maxpool_output_pipe_1021_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal sample_req, sample_ack : BooleanArray( 9 downto 0);
      signal update_req, update_ack : BooleanArray( 9 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 9 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1014_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_697_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_700_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_703_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_706_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_709_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_712_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_715_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_718_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1021_inst_req_0;
      WPIPE_maxpool_output_pipe_1014_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_697_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_700_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_703_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_706_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_709_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_712_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_715_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_718_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1021_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1014_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_697_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_700_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_703_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_706_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_709_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_712_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_715_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_718_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1021_inst_req_1;
      WPIPE_maxpool_output_pipe_1014_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_697_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_700_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_703_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_706_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_709_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_712_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_715_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_718_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1021_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      data_in <= tmp44x_xi_1013 & conv50_696 & conv44_686 & conv38_676 & conv32_666 & conv26_656 & conv20_646 & conv14_636 & conv8_626 & tmp49x_xi_1020;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 10, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 3,
      data_width => 8,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendModule is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
    output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendModule;
architecture sendModule_arch of sendModule is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendModule_CP_7437_start: Boolean;
  signal sendModule_CP_7437_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_output_pipe_2965_inst_req_1 : boolean;
  signal RPIPE_output_pipe_2965_inst_ack_1 : boolean;
  signal RPIPE_output_pipe_2971_inst_req_0 : boolean;
  signal RPIPE_output_pipe_2971_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_2971_inst_req_1 : boolean;
  signal array_obj_ref_3043_index_offset_ack_1 : boolean;
  signal RPIPE_output_pipe_2971_inst_ack_1 : boolean;
  signal phi_stmt_2991_req_0 : boolean;
  signal n_chl_3014_2990_buf_ack_1 : boolean;
  signal n_address_3027_2985_buf_req_1 : boolean;
  signal array_obj_ref_3043_index_offset_req_1 : boolean;
  signal phi_stmt_2981_req_1 : boolean;
  signal n_count_3035_2995_buf_req_0 : boolean;
  signal RPIPE_output_pipe_2968_inst_req_0 : boolean;
  signal RPIPE_output_pipe_2968_inst_ack_0 : boolean;
  signal phi_stmt_2986_req_1 : boolean;
  signal array_obj_ref_3043_index_offset_req_0 : boolean;
  signal n_count_3035_2995_buf_req_1 : boolean;
  signal n_chl_3014_2990_buf_req_0 : boolean;
  signal phi_stmt_2981_ack_0 : boolean;
  signal n_chl_3014_2990_buf_req_1 : boolean;
  signal n_count_3035_2995_buf_ack_0 : boolean;
  signal phi_stmt_2991_ack_0 : boolean;
  signal RPIPE_output_pipe_2965_inst_ack_0 : boolean;
  signal n_chl_3014_2990_buf_ack_0 : boolean;
  signal do_while_stmt_2979_branch_req_0 : boolean;
  signal RPIPE_output_pipe_2965_inst_req_0 : boolean;
  signal phi_stmt_2991_req_1 : boolean;
  signal phi_stmt_2986_ack_0 : boolean;
  signal SUB_u32_u32_3000_inst_ack_1 : boolean;
  signal n_count_3035_2995_buf_ack_1 : boolean;
  signal phi_stmt_2981_req_0 : boolean;
  signal addr_of_3044_final_reg_ack_1 : boolean;
  signal addr_of_3044_final_reg_req_1 : boolean;
  signal RPIPE_output_pipe_2968_inst_ack_1 : boolean;
  signal type_cast_3017_inst_ack_1 : boolean;
  signal type_cast_3017_inst_req_1 : boolean;
  signal RPIPE_output_pipe_2968_inst_req_1 : boolean;
  signal SUB_u32_u32_3000_inst_ack_0 : boolean;
  signal addr_of_3044_final_reg_ack_0 : boolean;
  signal addr_of_3044_final_reg_req_0 : boolean;
  signal type_cast_3017_inst_ack_0 : boolean;
  signal SUB_u32_u32_3000_inst_req_0 : boolean;
  signal type_cast_3017_inst_req_0 : boolean;
  signal SUB_u32_u32_3000_inst_req_1 : boolean;
  signal n_address_3027_2985_buf_ack_0 : boolean;
  signal phi_stmt_2986_req_0 : boolean;
  signal n_address_3027_2985_buf_req_0 : boolean;
  signal ptr_deref_3048_load_0_req_0 : boolean;
  signal ptr_deref_3048_load_0_ack_0 : boolean;
  signal array_obj_ref_3043_index_offset_ack_0 : boolean;
  signal n_address_3027_2985_buf_ack_1 : boolean;
  signal ptr_deref_3048_load_0_req_1 : boolean;
  signal ptr_deref_3048_load_0_ack_1 : boolean;
  signal RPIPE_output_pipe_3051_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3051_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3051_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3051_inst_ack_1 : boolean;
  signal slice_3055_inst_req_0 : boolean;
  signal slice_3055_inst_ack_0 : boolean;
  signal slice_3055_inst_req_1 : boolean;
  signal slice_3055_inst_ack_1 : boolean;
  signal slice_3059_inst_req_0 : boolean;
  signal slice_3059_inst_ack_0 : boolean;
  signal slice_3059_inst_req_1 : boolean;
  signal slice_3059_inst_ack_1 : boolean;
  signal slice_3063_inst_req_0 : boolean;
  signal slice_3063_inst_ack_0 : boolean;
  signal slice_3063_inst_req_1 : boolean;
  signal slice_3063_inst_ack_1 : boolean;
  signal slice_3067_inst_req_0 : boolean;
  signal slice_3067_inst_ack_0 : boolean;
  signal slice_3067_inst_req_1 : boolean;
  signal slice_3067_inst_ack_1 : boolean;
  signal EQ_u2_u1_3078_inst_req_0 : boolean;
  signal EQ_u2_u1_3078_inst_ack_0 : boolean;
  signal EQ_u2_u1_3078_inst_req_1 : boolean;
  signal EQ_u2_u1_3078_inst_ack_1 : boolean;
  signal W_output_data_2983_delayed_14_0_3080_inst_req_0 : boolean;
  signal W_output_data_2983_delayed_14_0_3080_inst_ack_0 : boolean;
  signal W_output_data_2983_delayed_14_0_3080_inst_req_1 : boolean;
  signal W_output_data_2983_delayed_14_0_3080_inst_ack_1 : boolean;
  signal EQ_u2_u1_3092_inst_req_0 : boolean;
  signal EQ_u2_u1_3092_inst_ack_0 : boolean;
  signal EQ_u2_u1_3092_inst_req_1 : boolean;
  signal EQ_u2_u1_3092_inst_ack_1 : boolean;
  signal W_output_data_2991_delayed_14_0_3094_inst_req_0 : boolean;
  signal W_output_data_2991_delayed_14_0_3094_inst_ack_0 : boolean;
  signal W_output_data_2991_delayed_14_0_3094_inst_req_1 : boolean;
  signal W_output_data_2991_delayed_14_0_3094_inst_ack_1 : boolean;
  signal EQ_u2_u1_3106_inst_req_0 : boolean;
  signal EQ_u2_u1_3106_inst_ack_0 : boolean;
  signal EQ_u2_u1_3106_inst_req_1 : boolean;
  signal EQ_u2_u1_3106_inst_ack_1 : boolean;
  signal W_output_data_2999_delayed_14_0_3108_inst_req_0 : boolean;
  signal W_output_data_2999_delayed_14_0_3108_inst_ack_0 : boolean;
  signal W_output_data_2999_delayed_14_0_3108_inst_req_1 : boolean;
  signal W_output_data_2999_delayed_14_0_3108_inst_ack_1 : boolean;
  signal EQ_u2_u1_3120_inst_req_0 : boolean;
  signal EQ_u2_u1_3120_inst_ack_0 : boolean;
  signal EQ_u2_u1_3120_inst_req_1 : boolean;
  signal EQ_u2_u1_3120_inst_ack_1 : boolean;
  signal W_output_data_3007_delayed_14_0_3122_inst_req_0 : boolean;
  signal W_output_data_3007_delayed_14_0_3122_inst_ack_0 : boolean;
  signal W_output_data_3007_delayed_14_0_3122_inst_req_1 : boolean;
  signal W_output_data_3007_delayed_14_0_3122_inst_ack_1 : boolean;
  signal W_fetch_addr_3011_delayed_8_0_3131_inst_req_0 : boolean;
  signal W_fetch_addr_3011_delayed_8_0_3131_inst_ack_0 : boolean;
  signal W_fetch_addr_3011_delayed_8_0_3131_inst_req_1 : boolean;
  signal W_fetch_addr_3011_delayed_8_0_3131_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3142_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3142_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3142_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3142_inst_ack_1 : boolean;
  signal ptr_deref_3135_store_0_req_0 : boolean;
  signal ptr_deref_3135_store_0_ack_0 : boolean;
  signal ptr_deref_3135_store_0_req_1 : boolean;
  signal ptr_deref_3135_store_0_ack_1 : boolean;
  signal SUB_u16_u16_3147_inst_req_0 : boolean;
  signal SUB_u16_u16_3147_inst_ack_0 : boolean;
  signal SUB_u16_u16_3147_inst_req_1 : boolean;
  signal SUB_u16_u16_3147_inst_ack_1 : boolean;
  signal do_while_stmt_2979_branch_ack_0 : boolean;
  signal do_while_stmt_2979_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3159_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3159_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3159_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3159_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendModule_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendModule_CP_7437_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendModule_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_7437_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendModule_CP_7437_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_7437_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendModule_CP_7437: Block -- control-path 
    signal sendModule_CP_7437_elements: BooleanArray(170 downto 0);
    -- 
  begin -- 
    sendModule_CP_7437_elements(0) <= sendModule_CP_7437_start;
    sendModule_CP_7437_symbol <= sendModule_CP_7437_elements(170);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2963/$entry
      -- CP-element group 0: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/$entry
      -- CP-element group 0: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978__entry__
      -- CP-element group 0: 	 branch_block_stmt_2963/branch_block_stmt_2963__entry__
      -- CP-element group 0: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_sample_start_
      -- 
    rr_7461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(0), ack => RPIPE_output_pipe_2965_inst_req_0); -- 
    -- CP-element group 1:  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	168 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	169 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2963/do_while_stmt_2979__exit__
      -- CP-element group 1: 	 branch_block_stmt_2963/assign_stmt_3161__entry__
      -- CP-element group 1: 	 branch_block_stmt_2963/assign_stmt_3161/$entry
      -- CP-element group 1: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Sample/req
      -- 
    req_8068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(1), ack => WPIPE_input_done_pipe_3159_inst_req_0); -- 
    sendModule_CP_7437_elements(1) <= sendModule_CP_7437_elements(168);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_sample_completed_
      -- 
    ra_7462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_2965_inst_ack_0, ack => sendModule_CP_7437_elements(2)); -- 
    cr_7466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(2), ack => RPIPE_output_pipe_2965_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2965_update_completed_
      -- 
    ca_7467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_2965_inst_ack_1, ack => sendModule_CP_7437_elements(3)); -- 
    rr_7475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(3), ack => RPIPE_output_pipe_2968_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Update/cr
      -- 
    ra_7476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_2968_inst_ack_0, ack => sendModule_CP_7437_elements(4)); -- 
    cr_7480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(4), ack => RPIPE_output_pipe_2968_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2968_Update/ca
      -- 
    ca_7481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_2968_inst_ack_1, ack => sendModule_CP_7437_elements(5)); -- 
    rr_7489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(5), ack => RPIPE_output_pipe_2971_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_sample_completed_
      -- 
    ra_7490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_2971_inst_ack_0, ack => sendModule_CP_7437_elements(6)); -- 
    cr_7494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(6), ack => RPIPE_output_pipe_2971_inst_req_1); -- 
    -- CP-element group 7:  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2963/do_while_stmt_2979__entry__
      -- CP-element group 7: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/$exit
      -- CP-element group 7: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978/RPIPE_output_pipe_2971_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2963/assign_stmt_2966_to_assign_stmt_2978__exit__
      -- 
    ca_7495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_2971_inst_ack_1, ack => sendModule_CP_7437_elements(7)); -- 
    -- CP-element group 8:  transition  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979__entry__
      -- CP-element group 8: 	 branch_block_stmt_2963/do_while_stmt_2979/$entry
      -- 
    sendModule_CP_7437_elements(8) <= sendModule_CP_7437_elements(7);
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	168 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979__exit__
      -- 
    -- Element group sendModule_CP_7437_elements(9) is bound as output of CP function.
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_back
      -- 
    -- Element group sendModule_CP_7437_elements(10) is bound as output of CP function.
    -- CP-element group 11:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	167 
    -- CP-element group 11: 	166 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_2963/do_while_stmt_2979/condition_done
      -- CP-element group 11: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_exit/$entry
      -- CP-element group 11: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_taken/$entry
      -- 
    sendModule_CP_7437_elements(11) <= sendModule_CP_7437_elements(16);
    -- CP-element group 12:  branch  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	165 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_body_done
      -- 
    sendModule_CP_7437_elements(12) <= sendModule_CP_7437_elements(165);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	25 
    -- CP-element group 13: 	44 
    -- CP-element group 13: 	63 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/back_edge_to_loop_body
      -- 
    sendModule_CP_7437_elements(13) <= sendModule_CP_7437_elements(10);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14: 	46 
    -- CP-element group 14: 	65 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/first_time_through_loop_body
      -- 
    sendModule_CP_7437_elements(14) <= sendModule_CP_7437_elements(8);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	85 
    -- CP-element group 15: 	80 
    -- CP-element group 15: 	95 
    -- CP-element group 15: 	76 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	159 
    -- CP-element group 15: 	163 
    -- CP-element group 15: 	86 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	39 
    -- CP-element group 15: 	57 
    -- CP-element group 15: 	58 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/loop_body_start
      -- CP-element group 15: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/$entry
      -- 
    -- Element group sendModule_CP_7437_elements(15) is bound as output of CP function.
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	79 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	162 
    -- CP-element group 16: 	163 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/condition_evaluated
      -- 
    condition_evaluated_7510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_7510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(16), ack => do_while_stmt_2979_branch_req_0); -- 
    sendModule_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(79) & sendModule_CP_7437_elements(20) & sendModule_CP_7437_elements(162) & sendModule_CP_7437_elements(163);
      gj_sendModule_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	38 
    -- CP-element group 17: 	57 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	59 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_sample_start__ps
      -- CP-element group 17: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/aggregated_phi_sample_req
      -- 
    sendModule_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(21) & sendModule_CP_7437_elements(38) & sendModule_CP_7437_elements(57) & sendModule_CP_7437_elements(20);
      gj_sendModule_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	23 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	60 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	81 
    -- CP-element group 18: 	77 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	57 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/aggregated_phi_sample_ack
      -- CP-element group 18: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_sample_completed_
      -- 
    sendModule_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(23) & sendModule_CP_7437_elements(41) & sendModule_CP_7437_elements(60);
      gj_sendModule_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	39 
    -- CP-element group 19: 	58 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	61 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_update_start__ps
      -- CP-element group 19: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/aggregated_phi_update_req
      -- 
    sendModule_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(22) & sendModule_CP_7437_elements(39) & sendModule_CP_7437_elements(58);
      gj_sendModule_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	62 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/aggregated_phi_update_ack
      -- 
    sendModule_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(24) & sendModule_CP_7437_elements(43) & sendModule_CP_7437_elements(62);
      gj_sendModule_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	83 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_sample_start_
      -- 
    sendModule_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(83) & sendModule_CP_7437_elements(79) & sendModule_CP_7437_elements(18);
      gj_sendModule_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	117 
    -- CP-element group 22: 	133 
    -- CP-element group 22: 	125 
    -- CP-element group 22: 	87 
    -- CP-element group 22: 	141 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	19 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_update_start_
      -- 
    sendModule_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(117) & sendModule_CP_7437_elements(133) & sendModule_CP_7437_elements(125) & sendModule_CP_7437_elements(87) & sendModule_CP_7437_elements(141);
      gj_sendModule_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	18 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7437_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	131 
    -- CP-element group 24: 	123 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	87 
    -- CP-element group 24: 	115 
    -- CP-element group 24: 	139 
    -- CP-element group 24:  members (15) 
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_resize_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_resize_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_resize_1/index_resize_req
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_scale_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_scale_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_resized_1
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_scaled_1
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_computed_1
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Sample/req
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_resize_1/index_resize_ack
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_scale_1/scale_rename_ack
      -- CP-element group 24: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_index_scale_1/scale_rename_req
      -- 
    req_7700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(24), ack => array_obj_ref_3043_index_offset_req_0); -- 
    -- Element group sendModule_CP_7437_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	13 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_loopback_trigger
      -- 
    sendModule_CP_7437_elements(25) <= sendModule_CP_7437_elements(13);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_loopback_sample_req
      -- CP-element group 26: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_loopback_sample_req_ps
      -- 
    phi_stmt_2981_loopback_sample_req_7525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2981_loopback_sample_req_7525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(26), ack => phi_stmt_2981_req_1); -- 
    -- Element group sendModule_CP_7437_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	14 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_entry_trigger
      -- 
    sendModule_CP_7437_elements(27) <= sendModule_CP_7437_elements(14);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_entry_sample_req_ps
      -- CP-element group 28: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_entry_sample_req
      -- 
    phi_stmt_2981_entry_sample_req_7528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2981_entry_sample_req_7528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(28), ack => phi_stmt_2981_req_0); -- 
    -- Element group sendModule_CP_7437_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_phi_mux_ack_ps
      -- CP-element group 29: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2981_phi_mux_ack
      -- 
    phi_stmt_2981_phi_mux_ack_7531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2981_ack_0, ack => sendModule_CP_7437_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_sample_start__ps
      -- 
    -- Element group sendModule_CP_7437_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_update_start_
      -- CP-element group 31: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_update_start__ps
      -- 
    -- Element group sendModule_CP_7437_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_update_completed__ps
      -- 
    sendModule_CP_7437_elements(32) <= sendModule_CP_7437_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2984_update_completed_
      -- 
    -- Element group sendModule_CP_7437_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => sendModule_CP_7437_elements(31), ack => sendModule_CP_7437_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Sample/req
      -- 
    req_7552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(34), ack => n_address_3027_2985_buf_req_0); -- 
    -- Element group sendModule_CP_7437_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Update/req
      -- CP-element group 35: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_update_start_
      -- CP-element group 35: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Update/$entry
      -- 
    req_7557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(35), ack => n_address_3027_2985_buf_req_1); -- 
    -- Element group sendModule_CP_7437_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Sample/ack
      -- 
    ack_7553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_3027_2985_buf_ack_0, ack => sendModule_CP_7437_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_address_2985_Update/ack
      -- 
    ack_7558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_3027_2985_buf_ack_1, ack => sendModule_CP_7437_elements(37)); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	79 
    -- CP-element group 38: 	18 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	17 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_sample_start_
      -- 
    sendModule_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(79) & sendModule_CP_7437_elements(18);
      gj_sendModule_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	15 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	43 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	19 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_update_start_
      -- 
    sendModule_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(43);
      gj_sendModule_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_sample_start__ps
      -- 
    sendModule_CP_7437_elements(40) <= sendModule_CP_7437_elements(17);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	18 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7437_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_update_start__ps
      -- 
    sendModule_CP_7437_elements(42) <= sendModule_CP_7437_elements(19);
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	39 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_update_completed__ps
      -- 
    -- Element group sendModule_CP_7437_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	13 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_loopback_trigger
      -- 
    sendModule_CP_7437_elements(44) <= sendModule_CP_7437_elements(13);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_loopback_sample_req_ps
      -- 
    phi_stmt_2986_loopback_sample_req_7569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2986_loopback_sample_req_7569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(45), ack => phi_stmt_2986_req_1); -- 
    -- Element group sendModule_CP_7437_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	14 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_entry_trigger
      -- 
    sendModule_CP_7437_elements(46) <= sendModule_CP_7437_elements(14);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_entry_sample_req_ps
      -- CP-element group 47: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_entry_sample_req
      -- 
    phi_stmt_2986_entry_sample_req_7572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2986_entry_sample_req_7572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(47), ack => phi_stmt_2986_req_0); -- 
    -- Element group sendModule_CP_7437_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_phi_mux_ack_ps
      -- CP-element group 48: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2986_phi_mux_ack
      -- 
    phi_stmt_2986_phi_mux_ack_7575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2986_ack_0, ack => sendModule_CP_7437_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_sample_start_
      -- 
    -- Element group sendModule_CP_7437_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_update_start_
      -- 
    -- Element group sendModule_CP_7437_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_update_completed__ps
      -- 
    sendModule_CP_7437_elements(51) <= sendModule_CP_7437_elements(52);
    -- CP-element group 52:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	51 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2989_update_completed_
      -- 
    -- Element group sendModule_CP_7437_elements(52) is a control-delay.
    cp_element_52_delay: control_delay_element  generic map(name => " 52_delay", delay_value => 1)  port map(req => sendModule_CP_7437_elements(50), ack => sendModule_CP_7437_elements(52), clk => clk, reset =>reset);
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Sample/req
      -- CP-element group 53: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_sample_start__ps
      -- 
    req_7596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(53), ack => n_chl_3014_2990_buf_req_0); -- 
    -- Element group sendModule_CP_7437_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_update_start_
      -- CP-element group 54: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Update/req
      -- CP-element group 54: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_update_start__ps
      -- CP-element group 54: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Update/$entry
      -- 
    req_7601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(54), ack => n_chl_3014_2990_buf_req_1); -- 
    -- Element group sendModule_CP_7437_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Sample/ack
      -- 
    ack_7597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3014_2990_buf_ack_0, ack => sendModule_CP_7437_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_chl_2990_Update/$exit
      -- 
    ack_7602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3014_2990_buf_ack_1, ack => sendModule_CP_7437_elements(56)); -- 
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	15 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	79 
    -- CP-element group 57: 	18 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	17 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_sample_start_
      -- 
    sendModule_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(79) & sendModule_CP_7437_elements(18);
      gj_sendModule_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	15 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	62 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	19 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_update_start_
      -- 
    sendModule_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(62);
      gj_sendModule_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	17 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_sample_start__ps
      -- 
    sendModule_CP_7437_elements(59) <= sendModule_CP_7437_elements(17);
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	18 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7437_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_update_start__ps
      -- 
    sendModule_CP_7437_elements(61) <= sendModule_CP_7437_elements(19);
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	20 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	58 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_update_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_update_completed_
      -- 
    -- Element group sendModule_CP_7437_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	13 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_loopback_trigger
      -- 
    sendModule_CP_7437_elements(63) <= sendModule_CP_7437_elements(13);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_loopback_sample_req_ps
      -- CP-element group 64: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_loopback_sample_req
      -- 
    phi_stmt_2991_loopback_sample_req_7613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2991_loopback_sample_req_7613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(64), ack => phi_stmt_2991_req_1); -- 
    -- Element group sendModule_CP_7437_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	14 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_entry_trigger
      -- 
    sendModule_CP_7437_elements(65) <= sendModule_CP_7437_elements(14);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_entry_sample_req
      -- CP-element group 66: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_entry_sample_req_ps
      -- 
    phi_stmt_2991_entry_sample_req_7616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2991_entry_sample_req_7616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(66), ack => phi_stmt_2991_req_0); -- 
    -- Element group sendModule_CP_7437_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_phi_mux_ack_ps
      -- CP-element group 67: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/phi_stmt_2991_phi_mux_ack
      -- 
    phi_stmt_2991_phi_mux_ack_7619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2991_ack_0, ack => sendModule_CP_7437_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_sample_start__ps
      -- 
    -- Element group sendModule_CP_7437_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_update_start__ps
      -- 
    -- Element group sendModule_CP_7437_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_update_completed__ps
      -- 
    sendModule_CP_7437_elements(70) <= sendModule_CP_7437_elements(71);
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	70 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_2994_update_completed_
      -- 
    -- Element group sendModule_CP_7437_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => sendModule_CP_7437_elements(69), ack => sendModule_CP_7437_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Sample/req
      -- 
    req_7640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(72), ack => n_count_3035_2995_buf_req_0); -- 
    -- Element group sendModule_CP_7437_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_update_start__ps
      -- CP-element group 73: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Update/req
      -- 
    req_7645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(73), ack => n_count_3035_2995_buf_req_1); -- 
    -- Element group sendModule_CP_7437_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Sample/ack
      -- 
    ack_7641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_3035_2995_buf_ack_0, ack => sendModule_CP_7437_elements(74)); -- 
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/R_n_count_2995_Update/ack
      -- 
    ack_7646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_3035_2995_buf_ack_1, ack => sendModule_CP_7437_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	15 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_sample_start_
      -- 
    rr_7655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(76), ack => SUB_u32_u32_3000_inst_req_0); -- 
    sendModule_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(78);
      gj_sendModule_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	18 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Update/cr
      -- 
    cr_7660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(77), ack => SUB_u32_u32_3000_inst_req_1); -- 
    sendModule_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(18) & sendModule_CP_7437_elements(79);
      gj_sendModule_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Sample/ra
      -- 
    ra_7656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3000_inst_ack_0, ack => sendModule_CP_7437_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	16 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	21 
    -- CP-element group 79: 	38 
    -- CP-element group 79: 	57 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u32_u32_3000_Update/ca
      -- 
    ca_7661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3000_inst_ack_1, ack => sendModule_CP_7437_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	15 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Sample/rr
      -- 
    rr_7669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(80), ack => type_cast_3017_inst_req_0); -- 
    sendModule_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(82);
      gj_sendModule_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	18 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_update_start_
      -- CP-element group 81: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Update/$entry
      -- 
    cr_7674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(81), ack => type_cast_3017_inst_req_1); -- 
    sendModule_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(18) & sendModule_CP_7437_elements(83);
      gj_sendModule_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Sample/ra
      -- 
    ra_7670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3017_inst_ack_0, ack => sendModule_CP_7437_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	165 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	21 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/type_cast_3017_Update/$exit
      -- 
    ca_7675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3017_inst_ack_1, ack => sendModule_CP_7437_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	88 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	89 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	89 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_request/req
      -- CP-element group 84: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_request/$entry
      -- 
    req_7715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(84), ack => addr_of_3044_final_reg_req_0); -- 
    sendModule_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(88) & sendModule_CP_7437_elements(89);
      gj_sendModule_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	15 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	93 
    -- CP-element group 85: 	149 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	90 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_complete/req
      -- CP-element group 85: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_complete/$entry
      -- 
    req_7720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(85), ack => addr_of_3044_final_reg_req_1); -- 
    sendModule_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(93) & sendModule_CP_7437_elements(149);
      gj_sendModule_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	15 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	89 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Update/req
      -- CP-element group 86: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_update_start
      -- 
    req_7705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(86), ack => array_obj_ref_3043_index_offset_req_1); -- 
    sendModule_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(89);
      gj_sendModule_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	24 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	165 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	22 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Sample/ack
      -- 
    ack_7701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3043_index_offset_ack_0, ack => sendModule_CP_7437_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	84 
    -- CP-element group 88:  members (8) 
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/array_obj_ref_3043_base_plus_offset/$exit
      -- 
    ack_7706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3043_index_offset_ack_1, ack => sendModule_CP_7437_elements(88)); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	84 
    -- CP-element group 89: successors 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	84 
    -- CP-element group 89: 	86 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_request/ack
      -- CP-element group 89: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_request/$exit
      -- 
    ack_7716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3044_final_reg_ack_0, ack => sendModule_CP_7437_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	85 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	147 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/addr_of_3044_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_word_addrgen/root_register_ack
      -- CP-element group 90: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_base_address_resized
      -- 
    ack_7721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3044_final_reg_ack_1, ack => sendModule_CP_7437_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	157 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/word_access_start/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/word_access_start/word_0/rr
      -- 
    rr_7754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(91), ack => ptr_deref_3048_load_0_req_0); -- 
    sendModule_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(90) & sendModule_CP_7437_elements(157);
      gj_sendModule_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	101 
    -- CP-element group 92: 	105 
    -- CP-element group 92: 	109 
    -- CP-element group 92: 	113 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/word_access_complete/word_0/cr
      -- 
    cr_7765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(92), ack => ptr_deref_3048_load_0_req_1); -- 
    sendModule_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(101) & sendModule_CP_7437_elements(105) & sendModule_CP_7437_elements(109) & sendModule_CP_7437_elements(113);
      gj_sendModule_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	164 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	85 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/word_access_start/word_0/$exit
      -- CP-element group 93: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/word_access_start/$exit
      -- CP-element group 93: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Sample/word_access_start/word_0/ra
      -- 
    ra_7755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3048_load_0_ack_0, ack => sendModule_CP_7437_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	99 
    -- CP-element group 94: 	107 
    -- CP-element group 94: 	103 
    -- CP-element group 94: 	111 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/word_access_complete/$exit
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/word_access_complete/word_0/$exit
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/word_access_complete/word_0/ca
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/ptr_deref_3048_Merge/$entry
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/ptr_deref_3048_Merge/$exit
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/ptr_deref_3048_Merge/merge_req
      -- CP-element group 94: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_Update/ptr_deref_3048_Merge/merge_ack
      -- 
    ca_7766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3048_load_0_ack_1, ack => sendModule_CP_7437_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	15 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	98 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Sample/rr
      -- 
    rr_7779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(95), ack => RPIPE_output_pipe_3051_inst_req_0); -- 
    sendModule_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(98);
      gj_sendModule_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	121 
    -- CP-element group 96: 	129 
    -- CP-element group 96: 	137 
    -- CP-element group 96: 	145 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_update_start_
      -- CP-element group 96: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Update/cr
      -- 
    cr_7784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(96), ack => RPIPE_output_pipe_3051_inst_req_1); -- 
    sendModule_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(97) & sendModule_CP_7437_elements(121) & sendModule_CP_7437_elements(129) & sendModule_CP_7437_elements(137) & sendModule_CP_7437_elements(145);
      gj_sendModule_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	96 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Sample/ra
      -- 
    ra_7780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3051_inst_ack_0, ack => sendModule_CP_7437_elements(97)); -- 
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	119 
    -- CP-element group 98: 	135 
    -- CP-element group 98: 	127 
    -- CP-element group 98: 	143 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	95 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/RPIPE_output_pipe_3051_Update/ca
      -- 
    ca_7785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3051_inst_ack_1, ack => sendModule_CP_7437_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	94 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Sample/rr
      -- 
    rr_7793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(99), ack => slice_3055_inst_req_0); -- 
    sendModule_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(94) & sendModule_CP_7437_elements(101);
      gj_sendModule_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	153 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Update/cr
      -- 
    cr_7798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(100), ack => slice_3055_inst_req_1); -- 
    sendModule_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	92 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Sample/ra
      -- 
    ra_7794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3055_inst_ack_0, ack => sendModule_CP_7437_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	151 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3055_Update/ca
      -- 
    ca_7799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3055_inst_ack_1, ack => sendModule_CP_7437_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	94 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	105 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Sample/rr
      -- 
    rr_7807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(103), ack => slice_3059_inst_req_0); -- 
    sendModule_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(94) & sendModule_CP_7437_elements(105);
      gj_sendModule_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	153 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Update/cr
      -- 
    cr_7812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(104), ack => slice_3059_inst_req_1); -- 
    sendModule_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: marked-successors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	92 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Sample/ra
      -- 
    ra_7808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3059_inst_ack_0, ack => sendModule_CP_7437_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	151 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3059_Update/ca
      -- 
    ca_7813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3059_inst_ack_1, ack => sendModule_CP_7437_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	94 
    -- CP-element group 107: marked-predecessors 
    -- CP-element group 107: 	109 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Sample/rr
      -- 
    rr_7821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(107), ack => slice_3063_inst_req_0); -- 
    sendModule_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(94) & sendModule_CP_7437_elements(109);
      gj_sendModule_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	153 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_update_start_
      -- CP-element group 108: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Update/cr
      -- 
    cr_7826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(108), ack => slice_3063_inst_req_1); -- 
    sendModule_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: marked-successors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	92 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Sample/ra
      -- 
    ra_7822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3063_inst_ack_0, ack => sendModule_CP_7437_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	151 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3063_Update/ca
      -- 
    ca_7827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3063_inst_ack_1, ack => sendModule_CP_7437_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	94 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Sample/rr
      -- 
    rr_7835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(111), ack => slice_3067_inst_req_0); -- 
    sendModule_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(94) & sendModule_CP_7437_elements(113);
      gj_sendModule_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	153 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_update_start_
      -- CP-element group 112: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Update/cr
      -- 
    cr_7840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(112), ack => slice_3067_inst_req_1); -- 
    sendModule_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	92 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Sample/ra
      -- 
    ra_7836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3067_inst_ack_0, ack => sendModule_CP_7437_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	151 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/slice_3067_Update/ca
      -- 
    ca_7841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3067_inst_ack_1, ack => sendModule_CP_7437_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	24 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Sample/rr
      -- 
    rr_7849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(115), ack => EQ_u2_u1_3078_inst_req_0); -- 
    sendModule_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(24) & sendModule_CP_7437_elements(117);
      gj_sendModule_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	153 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_update_start_
      -- CP-element group 116: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Update/cr
      -- 
    cr_7854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(116), ack => EQ_u2_u1_3078_inst_req_1); -- 
    sendModule_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	22 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Sample/ra
      -- 
    ra_7850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3078_inst_ack_0, ack => sendModule_CP_7437_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	151 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3078_Update/ca
      -- 
    ca_7855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3078_inst_ack_1, ack => sendModule_CP_7437_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	98 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Sample/req
      -- 
    req_7863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(119), ack => W_output_data_2983_delayed_14_0_3080_inst_req_0); -- 
    sendModule_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(98) & sendModule_CP_7437_elements(121);
      gj_sendModule_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	153 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_update_start_
      -- CP-element group 120: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Update/req
      -- 
    req_7868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(120), ack => W_output_data_2983_delayed_14_0_3080_inst_req_1); -- 
    sendModule_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	96 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Sample/ack
      -- 
    ack_7864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_2983_delayed_14_0_3080_inst_ack_0, ack => sendModule_CP_7437_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	151 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3082_Update/ack
      -- 
    ack_7869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_2983_delayed_14_0_3080_inst_ack_1, ack => sendModule_CP_7437_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	24 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Sample/rr
      -- 
    rr_7877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(123), ack => EQ_u2_u1_3092_inst_req_0); -- 
    sendModule_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(24) & sendModule_CP_7437_elements(125);
      gj_sendModule_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	153 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_update_start_
      -- CP-element group 124: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Update/cr
      -- 
    cr_7882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(124), ack => EQ_u2_u1_3092_inst_req_1); -- 
    sendModule_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	22 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Sample/ra
      -- 
    ra_7878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3092_inst_ack_0, ack => sendModule_CP_7437_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	151 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3092_Update/ca
      -- 
    ca_7883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3092_inst_ack_1, ack => sendModule_CP_7437_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	98 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Sample/req
      -- 
    req_7891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(127), ack => W_output_data_2991_delayed_14_0_3094_inst_req_0); -- 
    sendModule_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(98) & sendModule_CP_7437_elements(129);
      gj_sendModule_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	153 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_update_start_
      -- CP-element group 128: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Update/req
      -- 
    req_7896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(128), ack => W_output_data_2991_delayed_14_0_3094_inst_req_1); -- 
    sendModule_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	96 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Sample/ack
      -- 
    ack_7892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_2991_delayed_14_0_3094_inst_ack_0, ack => sendModule_CP_7437_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	151 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3096_Update/ack
      -- 
    ack_7897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_2991_delayed_14_0_3094_inst_ack_1, ack => sendModule_CP_7437_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	24 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Sample/rr
      -- 
    rr_7905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(131), ack => EQ_u2_u1_3106_inst_req_0); -- 
    sendModule_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(24) & sendModule_CP_7437_elements(133);
      gj_sendModule_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	153 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_update_start_
      -- CP-element group 132: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Update/cr
      -- 
    cr_7910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(132), ack => EQ_u2_u1_3106_inst_req_1); -- 
    sendModule_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: 	22 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Sample/ra
      -- 
    ra_7906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3106_inst_ack_0, ack => sendModule_CP_7437_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	151 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3106_Update/ca
      -- 
    ca_7911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3106_inst_ack_1, ack => sendModule_CP_7437_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	98 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Sample/req
      -- 
    req_7919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(135), ack => W_output_data_2999_delayed_14_0_3108_inst_req_0); -- 
    sendModule_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(98) & sendModule_CP_7437_elements(137);
      gj_sendModule_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	153 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_update_start_
      -- CP-element group 136: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Update/req
      -- 
    req_7924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(136), ack => W_output_data_2999_delayed_14_0_3108_inst_req_1); -- 
    sendModule_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: 	96 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Sample/ack
      -- 
    ack_7920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_2999_delayed_14_0_3108_inst_ack_0, ack => sendModule_CP_7437_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	151 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3110_Update/ack
      -- 
    ack_7925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_2999_delayed_14_0_3108_inst_ack_1, ack => sendModule_CP_7437_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	24 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Sample/rr
      -- 
    rr_7933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(139), ack => EQ_u2_u1_3120_inst_req_0); -- 
    sendModule_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(24) & sendModule_CP_7437_elements(141);
      gj_sendModule_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	153 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_update_start_
      -- CP-element group 140: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Update/cr
      -- 
    cr_7938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(140), ack => EQ_u2_u1_3120_inst_req_1); -- 
    sendModule_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	22 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Sample/ra
      -- 
    ra_7934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3120_inst_ack_0, ack => sendModule_CP_7437_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	151 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/EQ_u2_u1_3120_Update/ca
      -- 
    ca_7939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3120_inst_ack_1, ack => sendModule_CP_7437_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	98 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Sample/req
      -- 
    req_7947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(143), ack => W_output_data_3007_delayed_14_0_3122_inst_req_0); -- 
    sendModule_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(98) & sendModule_CP_7437_elements(145);
      gj_sendModule_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	153 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_update_start_
      -- CP-element group 144: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Update/req
      -- 
    req_7952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(144), ack => W_output_data_3007_delayed_14_0_3122_inst_req_1); -- 
    sendModule_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	96 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Sample/ack
      -- 
    ack_7948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_3007_delayed_14_0_3122_inst_ack_0, ack => sendModule_CP_7437_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	151 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3124_Update/ack
      -- 
    ack_7953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data_3007_delayed_14_0_3122_inst_ack_1, ack => sendModule_CP_7437_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	90 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Sample/req
      -- 
    req_7961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(147), ack => W_fetch_addr_3011_delayed_8_0_3131_inst_req_0); -- 
    sendModule_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(90) & sendModule_CP_7437_elements(149);
      gj_sendModule_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	157 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_update_start_
      -- CP-element group 148: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Update/req
      -- 
    req_7966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(148), ack => W_fetch_addr_3011_delayed_8_0_3131_inst_req_1); -- 
    sendModule_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(157);
      gj_sendModule_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	85 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Sample/ack
      -- 
    ack_7962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr_3011_delayed_8_0_3131_inst_ack_0, ack => sendModule_CP_7437_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	155 
    -- CP-element group 150:  members (19) 
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/assign_stmt_3133_Update/ack
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_address_calculated
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_word_address_calculated
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_root_address_calculated
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_address_resized
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_addr_resize/$entry
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_addr_resize/$exit
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_addr_resize/base_resize_req
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_addr_resize/base_resize_ack
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_plus_offset/$entry
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_plus_offset/$exit
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_plus_offset/sum_rename_req
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_base_plus_offset/sum_rename_ack
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_word_addrgen/$entry
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_word_addrgen/$exit
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_word_addrgen/root_register_req
      -- CP-element group 150: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_word_addrgen/root_register_ack
      -- 
    ack_7967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr_3011_delayed_8_0_3131_inst_ack_1, ack => sendModule_CP_7437_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	118 
    -- CP-element group 151: 	130 
    -- CP-element group 151: 	134 
    -- CP-element group 151: 	122 
    -- CP-element group 151: 	126 
    -- CP-element group 151: 	106 
    -- CP-element group 151: 	102 
    -- CP-element group 151: 	110 
    -- CP-element group 151: 	114 
    -- CP-element group 151: 	138 
    -- CP-element group 151: 	142 
    -- CP-element group 151: 	146 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Sample/rr
      -- 
    rr_7975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(151), ack => CONCAT_u32_u64_3142_inst_req_0); -- 
    sendModule_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(118) & sendModule_CP_7437_elements(130) & sendModule_CP_7437_elements(134) & sendModule_CP_7437_elements(122) & sendModule_CP_7437_elements(126) & sendModule_CP_7437_elements(106) & sendModule_CP_7437_elements(102) & sendModule_CP_7437_elements(110) & sendModule_CP_7437_elements(114) & sendModule_CP_7437_elements(138) & sendModule_CP_7437_elements(142) & sendModule_CP_7437_elements(146) & sendModule_CP_7437_elements(153);
      gj_sendModule_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	157 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_update_start_
      -- CP-element group 152: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Update/cr
      -- 
    cr_7980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(152), ack => CONCAT_u32_u64_3142_inst_req_1); -- 
    sendModule_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(157);
      gj_sendModule_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	120 
    -- CP-element group 153: 	132 
    -- CP-element group 153: 	136 
    -- CP-element group 153: 	100 
    -- CP-element group 153: 	124 
    -- CP-element group 153: 	128 
    -- CP-element group 153: 	108 
    -- CP-element group 153: 	104 
    -- CP-element group 153: 	112 
    -- CP-element group 153: 	116 
    -- CP-element group 153: 	140 
    -- CP-element group 153: 	144 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Sample/ra
      -- 
    ra_7976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3142_inst_ack_0, ack => sendModule_CP_7437_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/CONCAT_u32_u64_3142_Update/ca
      -- 
    ca_7981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3142_inst_ack_1, ack => sendModule_CP_7437_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: 	164 
    -- CP-element group 155: 	150 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/ptr_deref_3135_Split/$entry
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/ptr_deref_3135_Split/$exit
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/ptr_deref_3135_Split/split_req
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/ptr_deref_3135_Split/split_ack
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/word_access_start/word_0/rr
      -- 
    rr_8019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(155), ack => ptr_deref_3135_store_0_req_0); -- 
    sendModule_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(154) & sendModule_CP_7437_elements(164) & sendModule_CP_7437_elements(150) & sendModule_CP_7437_elements(157);
      gj_sendModule_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_update_start_
      -- CP-element group 156: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/word_access_complete/word_0/cr
      -- 
    cr_8030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(156), ack => ptr_deref_3135_store_0_req_1); -- 
    sendModule_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(158);
      gj_sendModule_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	165 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	91 
    -- CP-element group 157: 	155 
    -- CP-element group 157: 	148 
    -- CP-element group 157: 	152 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Sample/word_access_start/word_0/ra
      -- CP-element group 157: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ring_reenable_memory_space_0
      -- 
    ra_8020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3135_store_0_ack_0, ack => sendModule_CP_7437_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	165 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (5) 
      -- CP-element group 158: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3135_Update/word_access_complete/word_0/ca
      -- 
    ca_8031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3135_store_0_ack_1, ack => sendModule_CP_7437_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	15 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Sample/rr
      -- 
    rr_8039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(159), ack => SUB_u16_u16_3147_inst_req_0); -- 
    sendModule_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(15) & sendModule_CP_7437_elements(161);
      gj_sendModule_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_update_start_
      -- CP-element group 160: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Update/cr
      -- 
    cr_8044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(160), ack => SUB_u16_u16_3147_inst_req_1); -- 
    sendModule_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7437_elements(162);
      gj_sendModule_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Sample/ra
      -- 
    ra_8040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3147_inst_ack_0, ack => sendModule_CP_7437_elements(161)); -- 
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	16 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/SUB_u16_u16_3147_Update/ca
      -- 
    ca_8045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3147_inst_ack_1, ack => sendModule_CP_7437_elements(162)); -- 
    -- CP-element group 163:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	15 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	16 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group sendModule_CP_7437_elements(163) is a control-delay.
    cp_element_163_delay: control_delay_element  generic map(name => " 163_delay", delay_value => 1)  port map(req => sendModule_CP_7437_elements(15), ack => sendModule_CP_7437_elements(163), clk => clk, reset =>reset);
    -- CP-element group 164:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	93 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	155 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/ptr_deref_3048_ptr_deref_3135_delay
      -- 
    -- Element group sendModule_CP_7437_elements(164) is a control-delay.
    cp_element_164_delay: control_delay_element  generic map(name => " 164_delay", delay_value => 1)  port map(req => sendModule_CP_7437_elements(93), ack => sendModule_CP_7437_elements(164), clk => clk, reset =>reset);
    -- CP-element group 165:  join  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	83 
    -- CP-element group 165: 	157 
    -- CP-element group 165: 	158 
    -- CP-element group 165: 	87 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	12 
    -- CP-element group 165:  members (1) 
      -- CP-element group 165: 	 branch_block_stmt_2963/do_while_stmt_2979/do_while_stmt_2979_loop_body/$exit
      -- 
    sendModule_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7437_elements(83) & sendModule_CP_7437_elements(157) & sendModule_CP_7437_elements(158) & sendModule_CP_7437_elements(87);
      gj_sendModule_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7437_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	11 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_exit/$exit
      -- CP-element group 166: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_exit/ack
      -- 
    ack_8052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2979_branch_ack_0, ack => sendModule_CP_7437_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	11 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_taken/$exit
      -- CP-element group 167: 	 branch_block_stmt_2963/do_while_stmt_2979/loop_taken/ack
      -- 
    ack_8056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2979_branch_ack_1, ack => sendModule_CP_7437_elements(167)); -- 
    -- CP-element group 168:  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	9 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	1 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_2963/do_while_stmt_2979/$exit
      -- 
    sendModule_CP_7437_elements(168) <= sendModule_CP_7437_elements(9);
    -- CP-element group 169:  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	1 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (6) 
      -- CP-element group 169: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_update_start_
      -- CP-element group 169: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Update/req
      -- 
    ack_8069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3159_inst_ack_0, ack => sendModule_CP_7437_elements(169)); -- 
    req_8073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7437_elements(169), ack => WPIPE_input_done_pipe_3159_inst_req_1); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (8) 
      -- CP-element group 170: 	 branch_block_stmt_2963/assign_stmt_3161__exit__
      -- CP-element group 170: 	 branch_block_stmt_2963/$exit
      -- CP-element group 170: 	 branch_block_stmt_2963/branch_block_stmt_2963__exit__
      -- CP-element group 170: 	 $exit
      -- CP-element group 170: 	 branch_block_stmt_2963/assign_stmt_3161/$exit
      -- CP-element group 170: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_2963/assign_stmt_3161/WPIPE_input_done_pipe_3159_Update/ack
      -- 
    ack_8074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3159_inst_ack_1, ack => sendModule_CP_7437_elements(170)); -- 
    sendModule_do_while_stmt_2979_terminator_8057: loop_terminator -- 
      generic map (name => " sendModule_do_while_stmt_2979_terminator_8057", max_iterations_in_flight =>15) 
      port map(loop_body_exit => sendModule_CP_7437_elements(12),loop_continue => sendModule_CP_7437_elements(167),loop_terminate => sendModule_CP_7437_elements(166),loop_back => sendModule_CP_7437_elements(10),loop_exit => sendModule_CP_7437_elements(9),clk => clk, reset => reset); -- 
    phi_stmt_2981_phi_seq_7559_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7437_elements(27);
      sendModule_CP_7437_elements(30)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7437_elements(30);
      sendModule_CP_7437_elements(31)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7437_elements(32);
      sendModule_CP_7437_elements(28) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7437_elements(25);
      sendModule_CP_7437_elements(34)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7437_elements(36);
      sendModule_CP_7437_elements(35)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7437_elements(37);
      sendModule_CP_7437_elements(26) <= phi_mux_reqs(1);
      phi_stmt_2981_phi_seq_7559 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2981_phi_seq_7559") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7437_elements(17), 
          phi_sample_ack => sendModule_CP_7437_elements(23), 
          phi_update_req => sendModule_CP_7437_elements(19), 
          phi_update_ack => sendModule_CP_7437_elements(24), 
          phi_mux_ack => sendModule_CP_7437_elements(29), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2986_phi_seq_7603_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7437_elements(46);
      sendModule_CP_7437_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7437_elements(49);
      sendModule_CP_7437_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7437_elements(51);
      sendModule_CP_7437_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7437_elements(44);
      sendModule_CP_7437_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7437_elements(55);
      sendModule_CP_7437_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7437_elements(56);
      sendModule_CP_7437_elements(45) <= phi_mux_reqs(1);
      phi_stmt_2986_phi_seq_7603 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2986_phi_seq_7603") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7437_elements(40), 
          phi_sample_ack => sendModule_CP_7437_elements(41), 
          phi_update_req => sendModule_CP_7437_elements(42), 
          phi_update_ack => sendModule_CP_7437_elements(43), 
          phi_mux_ack => sendModule_CP_7437_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2991_phi_seq_7647_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7437_elements(65);
      sendModule_CP_7437_elements(68)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7437_elements(68);
      sendModule_CP_7437_elements(69)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7437_elements(70);
      sendModule_CP_7437_elements(66) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7437_elements(63);
      sendModule_CP_7437_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7437_elements(74);
      sendModule_CP_7437_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7437_elements(75);
      sendModule_CP_7437_elements(64) <= phi_mux_reqs(1);
      phi_stmt_2991_phi_seq_7647 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2991_phi_seq_7647") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7437_elements(59), 
          phi_sample_ack => sendModule_CP_7437_elements(60), 
          phi_update_req => sendModule_CP_7437_elements(61), 
          phi_update_ack => sendModule_CP_7437_elements(62), 
          phi_mux_ack => sendModule_CP_7437_elements(67), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_7511_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= sendModule_CP_7437_elements(13);
        preds(1)  <= sendModule_CP_7437_elements(14);
        entry_tmerge_7511 : transition_merge -- 
          generic map(name => " entry_tmerge_7511")
          port map (preds => preds, symbol_out => sendModule_CP_7437_elements(15));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_3011_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_3025_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3033_wire : std_logic_vector(31 downto 0);
    signal AND_u32_u32_3072_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3138_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3141_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_3142_wire : std_logic_vector(63 downto 0);
    signal EQ_u2_u1_2982_2982_delayed_14_0_3079 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2990_2990_delayed_14_0_3093 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2998_2998_delayed_14_0_3107 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3006_3006_delayed_14_0_3121 : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_3041_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_2976_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_3154_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_3025_3025_delayed_1_0_3148 : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_2911_2911_delayed_1_0_3001 : std_logic_vector(31 downto 0);
    signal ULT_u16_u1_3152_wire : std_logic_vector(0 downto 0);
    signal address_2981 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3043_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3043_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3043_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3043_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3043_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3043_root_address : std_logic_vector(13 downto 0);
    signal cb_2969 : std_logic_vector(15 downto 0);
    signal chl_2986 : std_logic_vector(15 downto 0);
    signal chl_change_3006 : std_logic_vector(0 downto 0);
    signal chl_out_2972 : std_logic_vector(15 downto 0);
    signal continue_flag_3156 : std_logic_vector(0 downto 0);
    signal count_2991 : std_logic_vector(31 downto 0);
    signal fetch_addr_3011_delayed_8_0_3133 : std_logic_vector(31 downto 0);
    signal fetch_addr_3045 : std_logic_vector(31 downto 0);
    signal fetch_val_3049 : std_logic_vector(63 downto 0);
    signal konst_2999_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3010_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3030_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3032_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3040_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3071_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3077_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3091_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3105_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3119_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3146_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3160_wire_constant : std_logic_vector(7 downto 0);
    signal location_3074 : std_logic_vector(1 downto 0);
    signal max_count_2978 : std_logic_vector(31 downto 0);
    signal n_address_3027 : std_logic_vector(31 downto 0);
    signal n_address_3027_2985_buffered : std_logic_vector(31 downto 0);
    signal n_chl_3014 : std_logic_vector(15 downto 0);
    signal n_chl_3014_2990_buffered : std_logic_vector(15 downto 0);
    signal n_count_3035 : std_logic_vector(31 downto 0);
    signal n_count_3035_2995_buffered : std_logic_vector(31 downto 0);
    signal output_data_2983_delayed_14_0_3082 : std_logic_vector(15 downto 0);
    signal output_data_2991_delayed_14_0_3096 : std_logic_vector(15 downto 0);
    signal output_data_2999_delayed_14_0_3110 : std_logic_vector(15 downto 0);
    signal output_data_3007_delayed_14_0_3124 : std_logic_vector(15 downto 0);
    signal output_data_3052 : std_logic_vector(15 downto 0);
    signal ptr_deref_3048_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3048_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3048_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3048_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3048_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3135_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3135_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3135_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3135_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3135_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3135_word_offset_0 : std_logic_vector(13 downto 0);
    signal rb_2966 : std_logic_vector(15 downto 0);
    signal type_cast_2928_2928_delayed_1_0_3018 : std_logic_vector(31 downto 0);
    signal type_cast_2984_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2989_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2994_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3022_wire : std_logic_vector(31 downto 0);
    signal type_cast_3042_resized : std_logic_vector(13 downto 0);
    signal type_cast_3042_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3042_wire : std_logic_vector(63 downto 0);
    signal w1_3056 : std_logic_vector(15 downto 0);
    signal w2_3060 : std_logic_vector(15 downto 0);
    signal w3_3064 : std_logic_vector(15 downto 0);
    signal w4_3068 : std_logic_vector(15 downto 0);
    signal wb1_3088 : std_logic_vector(15 downto 0);
    signal wb2_3102 : std_logic_vector(15 downto 0);
    signal wb3_3116 : std_logic_vector(15 downto 0);
    signal wb4_3130 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_3043_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3043_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3043_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3043_resized_base_address <= "00000000000000";
    konst_2999_wire_constant <= "00000000000000000000000000000001";
    konst_3010_wire_constant <= "0000000000000001";
    konst_3030_wire_constant <= "00000000000000000000000000000000";
    konst_3032_wire_constant <= "00000000000000000000000000000001";
    konst_3040_wire_constant <= "00000000000000000000000000000010";
    konst_3071_wire_constant <= "00000000000000000000000000000011";
    konst_3077_wire_constant <= "00";
    konst_3091_wire_constant <= "01";
    konst_3105_wire_constant <= "10";
    konst_3119_wire_constant <= "11";
    konst_3146_wire_constant <= "0000000000000001";
    konst_3160_wire_constant <= "00000001";
    ptr_deref_3048_word_offset_0 <= "00000000000000";
    ptr_deref_3135_word_offset_0 <= "00000000000000";
    type_cast_2984_wire_constant <= "00000000000000000000000000000000";
    type_cast_2989_wire_constant <= "0000000000000000";
    type_cast_2994_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_2981: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2984_wire_constant & n_address_3027_2985_buffered;
      req <= phi_stmt_2981_req_0 & phi_stmt_2981_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2981",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2981_ack_0,
          idata => idata,
          odata => address_2981,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2981
    phi_stmt_2986: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2989_wire_constant & n_chl_3014_2990_buffered;
      req <= phi_stmt_2986_req_0 & phi_stmt_2986_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2986",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2986_ack_0,
          idata => idata,
          odata => chl_2986,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2986
    phi_stmt_2991: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2994_wire_constant & n_count_3035_2995_buffered;
      req <= phi_stmt_2991_req_0 & phi_stmt_2991_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2991",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2991_ack_0,
          idata => idata,
          odata => count_2991,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2991
    -- flow-through select operator MUX_3013_inst
    n_chl_3014 <= ADD_u16_u16_3011_wire when (chl_change_3006(0) /=  '0') else chl_2986;
    -- flow-through select operator MUX_3026_inst
    n_address_3027 <= type_cast_3022_wire when (chl_change_3006(0) /=  '0') else ADD_u32_u32_3025_wire;
    -- flow-through select operator MUX_3034_inst
    n_count_3035 <= konst_3030_wire_constant when (chl_change_3006(0) /=  '0') else ADD_u32_u32_3033_wire;
    -- flow-through select operator MUX_3087_inst
    wb1_3088 <= output_data_2983_delayed_14_0_3082 when (EQ_u2_u1_2982_2982_delayed_14_0_3079(0) /=  '0') else w1_3056;
    -- flow-through select operator MUX_3101_inst
    wb2_3102 <= output_data_2991_delayed_14_0_3096 when (EQ_u2_u1_2990_2990_delayed_14_0_3093(0) /=  '0') else w2_3060;
    -- flow-through select operator MUX_3115_inst
    wb3_3116 <= output_data_2999_delayed_14_0_3110 when (EQ_u2_u1_2998_2998_delayed_14_0_3107(0) /=  '0') else w3_3064;
    -- flow-through select operator MUX_3129_inst
    wb4_3130 <= output_data_3007_delayed_14_0_3124 when (EQ_u2_u1_3006_3006_delayed_14_0_3121(0) /=  '0') else w4_3068;
    slice_3055_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3055_inst_req_0;
      slice_3055_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3055_inst_req_1;
      slice_3055_inst_ack_1<= update_ack(0);
      slice_3055_inst: SliceSplitProtocol generic map(name => "slice_3055_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val_3049, dout => w1_3056, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3059_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3059_inst_req_0;
      slice_3059_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3059_inst_req_1;
      slice_3059_inst_ack_1<= update_ack(0);
      slice_3059_inst: SliceSplitProtocol generic map(name => "slice_3059_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val_3049, dout => w2_3060, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3063_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3063_inst_req_0;
      slice_3063_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3063_inst_req_1;
      slice_3063_inst_ack_1<= update_ack(0);
      slice_3063_inst: SliceSplitProtocol generic map(name => "slice_3063_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val_3049, dout => w3_3064, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3067_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3067_inst_req_0;
      slice_3067_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3067_inst_req_1;
      slice_3067_inst_ack_1<= update_ack(0);
      slice_3067_inst: SliceSplitProtocol generic map(name => "slice_3067_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val_3049, dout => w4_3068, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_fetch_addr_3011_delayed_8_0_3131_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr_3011_delayed_8_0_3131_inst_req_0;
      W_fetch_addr_3011_delayed_8_0_3131_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr_3011_delayed_8_0_3131_inst_req_1;
      W_fetch_addr_3011_delayed_8_0_3131_inst_ack_1<= rack(0);
      W_fetch_addr_3011_delayed_8_0_3131_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr_3011_delayed_8_0_3131_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr_3045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_3011_delayed_8_0_3133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data_2983_delayed_14_0_3080_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data_2983_delayed_14_0_3080_inst_req_0;
      W_output_data_2983_delayed_14_0_3080_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data_2983_delayed_14_0_3080_inst_req_1;
      W_output_data_2983_delayed_14_0_3080_inst_ack_1<= rack(0);
      W_output_data_2983_delayed_14_0_3080_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data_2983_delayed_14_0_3080_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data_3052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data_2983_delayed_14_0_3082,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data_2991_delayed_14_0_3094_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data_2991_delayed_14_0_3094_inst_req_0;
      W_output_data_2991_delayed_14_0_3094_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data_2991_delayed_14_0_3094_inst_req_1;
      W_output_data_2991_delayed_14_0_3094_inst_ack_1<= rack(0);
      W_output_data_2991_delayed_14_0_3094_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data_2991_delayed_14_0_3094_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data_3052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data_2991_delayed_14_0_3096,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data_2999_delayed_14_0_3108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data_2999_delayed_14_0_3108_inst_req_0;
      W_output_data_2999_delayed_14_0_3108_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data_2999_delayed_14_0_3108_inst_req_1;
      W_output_data_2999_delayed_14_0_3108_inst_ack_1<= rack(0);
      W_output_data_2999_delayed_14_0_3108_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data_2999_delayed_14_0_3108_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data_3052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data_2999_delayed_14_0_3110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data_3007_delayed_14_0_3122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data_3007_delayed_14_0_3122_inst_req_0;
      W_output_data_3007_delayed_14_0_3122_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data_3007_delayed_14_0_3122_inst_req_1;
      W_output_data_3007_delayed_14_0_3122_inst_ack_1<= rack(0);
      W_output_data_3007_delayed_14_0_3122_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data_3007_delayed_14_0_3122_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data_3052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data_3007_delayed_14_0_3124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3044_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3044_final_reg_req_0;
      addr_of_3044_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3044_final_reg_req_1;
      addr_of_3044_final_reg_ack_1<= rack(0);
      addr_of_3044_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3044_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3043_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_3045,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_3027_2985_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_3027_2985_buf_req_0;
      n_address_3027_2985_buf_ack_0<= wack(0);
      rreq(0) <= n_address_3027_2985_buf_req_1;
      n_address_3027_2985_buf_ack_1<= rack(0);
      n_address_3027_2985_buf : InterlockBuffer generic map ( -- 
        name => "n_address_3027_2985_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_3027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_3027_2985_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_3014_2990_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_3014_2990_buf_req_0;
      n_chl_3014_2990_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_3014_2990_buf_req_1;
      n_chl_3014_2990_buf_ack_1<= rack(0);
      n_chl_3014_2990_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_3014_2990_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_3014,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_3014_2990_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_count_3035_2995_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_3035_2995_buf_req_0;
      n_count_3035_2995_buf_ack_0<= wack(0);
      rreq(0) <= n_count_3035_2995_buf_req_1;
      n_count_3035_2995_buf_ack_1<= rack(0);
      n_count_3035_2995_buf : InterlockBuffer generic map ( -- 
        name => "n_count_3035_2995_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_3035,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_3035_2995_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2977_inst
    process(MUL_u16_u16_2976_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_2976_wire(15 downto 0);
      max_count_2978 <= tmp_var; -- 
    end process;
    type_cast_3017_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3017_inst_req_0;
      type_cast_3017_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3017_inst_req_1;
      type_cast_3017_inst_ack_1<= rack(0);
      type_cast_3017_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3017_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_2972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2928_2928_delayed_1_0_3018,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3022_inst
    process(n_chl_3014) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3014(15 downto 0);
      type_cast_3022_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3042_inst
    process(LSHR_u32_u32_3041_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3041_wire(31 downto 0);
      type_cast_3042_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3073_inst
    process(AND_u32_u32_3072_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := AND_u32_u32_3072_wire(1 downto 0);
      location_3074 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_3043_index_1_rename
    process(type_cast_3042_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3042_resized;
      ov(13 downto 0) := iv;
      type_cast_3042_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3043_index_1_resize
    process(type_cast_3042_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3042_wire;
      ov := iv(13 downto 0);
      type_cast_3042_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3043_root_address_inst
    process(array_obj_ref_3043_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3043_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3043_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3048_addr_0
    process(ptr_deref_3048_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3048_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3048_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3048_base_resize
    process(fetch_addr_3045) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_3045;
      ov := iv(13 downto 0);
      ptr_deref_3048_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3048_gather_scatter
    process(ptr_deref_3048_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3048_data_0;
      ov(63 downto 0) := iv;
      fetch_val_3049 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3048_root_address_inst
    process(ptr_deref_3048_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3048_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3048_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3135_addr_0
    process(ptr_deref_3135_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3135_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3135_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3135_base_resize
    process(fetch_addr_3011_delayed_8_0_3133) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_3011_delayed_8_0_3133;
      ov := iv(13 downto 0);
      ptr_deref_3135_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3135_gather_scatter
    process(CONCAT_u32_u64_3142_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3142_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3135_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3135_root_address_inst
    process(ptr_deref_3135_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3135_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3135_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_2979_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_3156;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2979_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2979_branch_req_0,
          ack0 => do_while_stmt_2979_branch_ack_0,
          ack1 => do_while_stmt_2979_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3011_inst
    process(chl_2986) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_2986, konst_3010_wire_constant, tmp_var);
      ADD_u16_u16_3011_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3025_inst
    process(address_2981, type_cast_2928_2928_delayed_1_0_3018) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_2981, type_cast_2928_2928_delayed_1_0_3018, tmp_var);
      ADD_u32_u32_3025_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3033_inst
    process(count_2991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_2991, konst_3032_wire_constant, tmp_var);
      ADD_u32_u32_3033_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_3072_inst
    process(address_2981) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address_2981, konst_3071_wire_constant, tmp_var);
      AND_u32_u32_3072_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3138_inst
    process(wb1_3088, wb2_3102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb1_3088, wb2_3102, tmp_var);
      CONCAT_u16_u32_3138_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3141_inst
    process(wb3_3116, wb4_3130) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb3_3116, wb4_3130, tmp_var);
      CONCAT_u16_u32_3141_wire <= tmp_var; --
    end process;
    -- shared split operator group (6) : CONCAT_u32_u64_3142_inst 
    ApConcat_group_6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3138_wire & CONCAT_u16_u32_3141_wire;
      CONCAT_u32_u64_3142_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3142_inst_req_0;
      CONCAT_u32_u64_3142_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3142_inst_req_1;
      CONCAT_u32_u64_3142_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_6_gI: SplitGuardInterface generic map(name => "ApConcat_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u2_u1_3078_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location_3074;
      EQ_u2_u1_2982_2982_delayed_14_0_3079 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3078_inst_req_0;
      EQ_u2_u1_3078_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3078_inst_req_1;
      EQ_u2_u1_3078_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : EQ_u2_u1_3092_inst 
    ApIntEq_group_8: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location_3074;
      EQ_u2_u1_2990_2990_delayed_14_0_3093 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3092_inst_req_0;
      EQ_u2_u1_3092_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3092_inst_req_1;
      EQ_u2_u1_3092_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_8_gI: SplitGuardInterface generic map(name => "ApIntEq_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : EQ_u2_u1_3106_inst 
    ApIntEq_group_9: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location_3074;
      EQ_u2_u1_2998_2998_delayed_14_0_3107 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3106_inst_req_0;
      EQ_u2_u1_3106_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3106_inst_req_1;
      EQ_u2_u1_3106_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_9_gI: SplitGuardInterface generic map(name => "ApIntEq_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : EQ_u2_u1_3120_inst 
    ApIntEq_group_10: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location_3074;
      EQ_u2_u1_3006_3006_delayed_14_0_3121 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3120_inst_req_0;
      EQ_u2_u1_3120_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3120_inst_req_1;
      EQ_u2_u1_3120_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_10_gI: SplitGuardInterface generic map(name => "ApIntEq_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- binary operator EQ_u32_u1_3005_inst
    process(count_2991, SUB_u32_u32_2911_2911_delayed_1_0_3001) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_2991, SUB_u32_u32_2911_2911_delayed_1_0_3001, tmp_var);
      chl_change_3006 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3041_inst
    process(address_2981) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address_2981, konst_3040_wire_constant, tmp_var);
      LSHR_u32_u32_3041_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2976_inst
    process(rb_2966, cb_2969) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(rb_2966, cb_2969, tmp_var);
      MUL_u16_u16_2976_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3154_inst
    process(chl_change_3006) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", chl_change_3006, tmp_var);
      NOT_u1_u1_3154_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_3155_inst
    process(ULT_u16_u1_3152_wire, NOT_u1_u1_3154_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ULT_u16_u1_3152_wire, NOT_u1_u1_3154_wire, tmp_var);
      continue_flag_3156 <= tmp_var; --
    end process;
    -- shared split operator group (16) : SUB_u16_u16_3147_inst 
    ApIntSub_group_16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= chl_out_2972;
      SUB_u16_u16_3025_3025_delayed_1_0_3148 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3147_inst_req_0;
      SUB_u16_u16_3147_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3147_inst_req_1;
      SUB_u16_u16_3147_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_16_gI: SplitGuardInterface generic map(name => "ApIntSub_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : SUB_u32_u32_3000_inst 
    ApIntSub_group_17: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= max_count_2978;
      SUB_u32_u32_2911_2911_delayed_1_0_3001 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3000_inst_req_0;
      SUB_u32_u32_3000_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3000_inst_req_1;
      SUB_u32_u32_3000_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_17_gI: SplitGuardInterface generic map(name => "ApIntSub_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- binary operator ULT_u16_u1_3152_inst
    process(chl_2986, SUB_u16_u16_3025_3025_delayed_1_0_3148) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(chl_2986, SUB_u16_u16_3025_3025_delayed_1_0_3148, tmp_var);
      ULT_u16_u1_3152_wire <= tmp_var; --
    end process;
    -- shared split operator group (19) : array_obj_ref_3043_index_offset 
    ApIntAdd_group_19: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3042_scaled;
      array_obj_ref_3043_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3043_index_offset_req_0;
      array_obj_ref_3043_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3043_index_offset_req_1;
      array_obj_ref_3043_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_19_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared load operator group (0) : ptr_deref_3048_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3048_load_0_req_0;
      ptr_deref_3048_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3048_load_0_req_1;
      ptr_deref_3048_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3048_word_address_0;
      ptr_deref_3048_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3135_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3135_store_0_req_0;
      ptr_deref_3135_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3135_store_0_req_1;
      ptr_deref_3135_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3135_word_address_0;
      data_in <= ptr_deref_3135_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_output_pipe_2971_inst RPIPE_output_pipe_2968_inst RPIPE_output_pipe_2965_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(47 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 2 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= RPIPE_output_pipe_2971_inst_req_0;
      reqL_unguarded(1) <= RPIPE_output_pipe_2968_inst_req_0;
      reqL_unguarded(0) <= RPIPE_output_pipe_2965_inst_req_0;
      RPIPE_output_pipe_2971_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_output_pipe_2968_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_output_pipe_2965_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= RPIPE_output_pipe_2971_inst_req_1;
      reqR_unguarded(1) <= RPIPE_output_pipe_2968_inst_req_1;
      reqR_unguarded(0) <= RPIPE_output_pipe_2965_inst_req_1;
      RPIPE_output_pipe_2971_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_output_pipe_2968_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_output_pipe_2965_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      chl_out_2972 <= data_out(47 downto 32);
      cb_2969 <= data_out(31 downto 16);
      rb_2966 <= data_out(15 downto 0);
      output_pipe_read_0_gI: SplitGuardInterface generic map(name => "output_pipe_read_0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_0: InputPortRevised -- 
        generic map ( name => "output_pipe_read_0", data_width => 16,  num_reqs => 3,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(1),
          oack => output_pipe_pipe_read_ack(1),
          odata => output_pipe_pipe_read_data(31 downto 16),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_output_pipe_3051_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_output_pipe_3051_inst_req_0;
      RPIPE_output_pipe_3051_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_output_pipe_3051_inst_req_1;
      RPIPE_output_pipe_3051_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      output_data_3052 <= data_out(15 downto 0);
      output_pipe_read_1_gI: SplitGuardInterface generic map(name => "output_pipe_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_1: InputPortRevised -- 
        generic map ( name => "output_pipe_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(0),
          oack => output_pipe_pipe_read_ack(0),
          odata => output_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3159_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3159_inst_req_0;
      WPIPE_input_done_pipe_3159_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3159_inst_req_1;
      WPIPE_input_done_pipe_3159_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3160_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendModule_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_1275_start: Boolean;
  signal timer_CP_1275_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_383_inst_req_0 : boolean;
  signal WPIPE_timer_req_383_inst_ack_0 : boolean;
  signal WPIPE_timer_req_383_inst_req_1 : boolean;
  signal WPIPE_timer_req_383_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_388_inst_req_0 : boolean;
  signal RPIPE_timer_resp_388_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_388_inst_req_1 : boolean;
  signal RPIPE_timer_resp_388_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_1275_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1275_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_1275_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1275_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_1275: Block -- control-path 
    signal timer_CP_1275_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_1275_elements(0) <= timer_CP_1275_start;
    timer_CP_1275_symbol <= timer_CP_1275_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_389/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_sample_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Sample/req
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_sample_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Sample/rr
      -- 
    rr_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(0), ack => RPIPE_timer_resp_388_inst_req_0); -- 
    req_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(0), ack => WPIPE_timer_req_383_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_sample_completed_
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_update_start_
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Sample/ack
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Update/$entry
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Update/req
      -- 
    ack_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_383_inst_ack_0, ack => timer_CP_1275_elements(1)); -- 
    req_1293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(1), ack => WPIPE_timer_req_383_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_update_completed_
      -- CP-element group 2: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Update/$exit
      -- CP-element group 2: 	 assign_stmt_386_to_assign_stmt_389/WPIPE_timer_req_383_Update/ack
      -- 
    ack_1294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_383_inst_ack_1, ack => timer_CP_1275_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_sample_completed_
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_update_start_
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Sample/ra
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Update/$entry
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Update/cr
      -- 
    ra_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_388_inst_ack_0, ack => timer_CP_1275_elements(3)); -- 
    cr_1307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(3), ack => RPIPE_timer_resp_388_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_update_completed_
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Update/$exit
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_389/RPIPE_timer_resp_388_Update/ca
      -- 
    ca_1308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_388_inst_ack_1, ack => timer_CP_1275_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_386_to_assign_stmt_389/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_1275_elements(2) & timer_CP_1275_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_1275_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_385_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_385_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_388_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_388_inst_req_0;
      RPIPE_timer_resp_388_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_388_inst_req_1;
      RPIPE_timer_resp_388_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_383_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_383_inst_req_0;
      WPIPE_timer_req_383_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_383_inst_req_1;
      WPIPE_timer_req_383_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_385_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_8970_start: Boolean;
  signal timerDaemon_CP_8970_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_3437_branch_req_0 : boolean;
  signal RPIPE_timer_req_3446_inst_ack_0 : boolean;
  signal RPIPE_timer_req_3446_inst_req_0 : boolean;
  signal do_while_stmt_3437_branch_ack_1 : boolean;
  signal do_while_stmt_3437_branch_ack_0 : boolean;
  signal WPIPE_timer_resp_3454_inst_ack_0 : boolean;
  signal nCOUNTER_3452_3443_buf_ack_0 : boolean;
  signal nCOUNTER_3452_3443_buf_req_0 : boolean;
  signal phi_stmt_3439_req_0 : boolean;
  signal RPIPE_timer_req_3446_inst_ack_1 : boolean;
  signal RPIPE_timer_req_3446_inst_req_1 : boolean;
  signal nCOUNTER_3452_3443_buf_ack_1 : boolean;
  signal nCOUNTER_3452_3443_buf_req_1 : boolean;
  signal phi_stmt_3439_req_1 : boolean;
  signal WPIPE_timer_resp_3454_inst_req_0 : boolean;
  signal phi_stmt_3439_ack_0 : boolean;
  signal WPIPE_timer_resp_3454_inst_req_1 : boolean;
  signal WPIPE_timer_resp_3454_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_8970_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_8970_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_8970_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_8970_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_8970: Block -- control-path 
    signal timerDaemon_CP_8970_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_8970_elements(0) <= timerDaemon_CP_8970_start;
    timerDaemon_CP_8970_symbol <= timerDaemon_CP_8970_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_3436/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3436/do_while_stmt_3437__entry__
      -- CP-element group 0: 	 branch_block_stmt_3436/branch_block_stmt_3436__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_3436/$exit
      -- CP-element group 1: 	 branch_block_stmt_3436/branch_block_stmt_3436__exit__
      -- CP-element group 1: 	 branch_block_stmt_3436/do_while_stmt_3437__exit__
      -- 
    timerDaemon_CP_8970_elements(1) <= timerDaemon_CP_8970_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_3436/do_while_stmt_3437/$entry
      -- CP-element group 2: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437__entry__
      -- 
    timerDaemon_CP_8970_elements(2) <= timerDaemon_CP_8970_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437__exit__
      -- 
    -- Element group timerDaemon_CP_8970_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_back
      -- 
    -- Element group timerDaemon_CP_8970_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_3436/do_while_stmt_3437/condition_done
      -- CP-element group 5: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_exit/$entry
      -- 
    timerDaemon_CP_8970_elements(5) <= timerDaemon_CP_8970_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_body_done
      -- 
    timerDaemon_CP_8970_elements(6) <= timerDaemon_CP_8970_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_8970_elements(7) <= timerDaemon_CP_8970_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_8970_elements(8) <= timerDaemon_CP_8970_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3444_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/$entry
      -- 
    -- Element group timerDaemon_CP_8970_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/condition_evaluated
      -- 
    condition_evaluated_8994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_8994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(10), ack => do_while_stmt_3437_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(14) & timerDaemon_CP_8970_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(9) & timerDaemon_CP_8970_elements(15) & timerDaemon_CP_8970_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3444_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(17) & timerDaemon_CP_8970_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(16) & timerDaemon_CP_8970_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(18) & timerDaemon_CP_8970_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(9) & timerDaemon_CP_8970_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(9) & timerDaemon_CP_8970_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_8970_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_8970_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_loopback_trigger
      -- 
    timerDaemon_CP_8970_elements(19) <= timerDaemon_CP_8970_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_loopback_sample_req
      -- 
    phi_stmt_3439_loopback_sample_req_9009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3439_loopback_sample_req_9009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(20), ack => phi_stmt_3439_req_1); -- 
    -- Element group timerDaemon_CP_8970_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_entry_trigger
      -- 
    timerDaemon_CP_8970_elements(21) <= timerDaemon_CP_8970_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_entry_sample_req
      -- 
    phi_stmt_3439_entry_sample_req_9012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3439_entry_sample_req_9012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(22), ack => phi_stmt_3439_req_0); -- 
    -- Element group timerDaemon_CP_8970_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3439_phi_mux_ack
      -- 
    phi_stmt_3439_phi_mux_ack_9015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3439_ack_0, ack => timerDaemon_CP_8970_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_sample_start_
      -- 
    -- Element group timerDaemon_CP_8970_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_update_start_
      -- 
    -- Element group timerDaemon_CP_8970_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_update_completed__ps
      -- 
    timerDaemon_CP_8970_elements(26) <= timerDaemon_CP_8970_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/type_cast_3442_update_completed_
      -- 
    -- Element group timerDaemon_CP_8970_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_8970_elements(25), ack => timerDaemon_CP_8970_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_sample_start__ps
      -- 
    req_9036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(28), ack => nCOUNTER_3452_3443_buf_req_0); -- 
    -- Element group timerDaemon_CP_8970_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_update_start_
      -- CP-element group 29: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Update/req
      -- CP-element group 29: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_update_start__ps
      -- 
    req_9041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(29), ack => nCOUNTER_3452_3443_buf_req_1); -- 
    -- Element group timerDaemon_CP_8970_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_sample_completed__ps
      -- 
    ack_9037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3452_3443_buf_ack_0, ack => timerDaemon_CP_8970_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/R_nCOUNTER_3443_update_completed__ps
      -- 
    ack_9042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3452_3443_buf_ack_1, ack => timerDaemon_CP_8970_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3444_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(9) & timerDaemon_CP_8970_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_sample_start_
      -- 
    rr_9055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(33), ack => RPIPE_timer_req_3446_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(11) & timerDaemon_CP_8970_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_update_start_
      -- CP-element group 34: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Update/$entry
      -- 
    cr_9060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(34), ack => RPIPE_timer_req_3446_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(13) & timerDaemon_CP_8970_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_sample_completed_
      -- 
    ra_9056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3446_inst_ack_0, ack => timerDaemon_CP_8970_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/RPIPE_timer_req_3446_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/phi_stmt_3444_update_completed_
      -- 
    ca_9061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3446_inst_ack_1, ack => timerDaemon_CP_8970_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Sample/req
      -- 
    req_9069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(37), ack => WPIPE_timer_resp_3454_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(18) & timerDaemon_CP_8970_elements(36) & timerDaemon_CP_8970_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_update_start_
      -- CP-element group 38: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Update/req
      -- 
    ack_9070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3454_inst_ack_0, ack => timerDaemon_CP_8970_elements(38)); -- 
    req_9074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_8970_elements(38), ack => WPIPE_timer_resp_3454_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/WPIPE_timer_resp_3454_Update/$exit
      -- 
    ack_9075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3454_inst_ack_1, ack => timerDaemon_CP_8970_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_8970_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_8970_elements(9), ack => timerDaemon_CP_8970_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3436/do_while_stmt_3437/do_while_stmt_3437_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_8970_elements(12) & timerDaemon_CP_8970_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_8970_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_exit/ack
      -- CP-element group 42: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_exit/$exit
      -- 
    ack_9080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3437_branch_ack_0, ack => timerDaemon_CP_8970_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_taken/ack
      -- CP-element group 43: 	 branch_block_stmt_3436/do_while_stmt_3437/loop_taken/$exit
      -- 
    ack_9084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3437_branch_ack_1, ack => timerDaemon_CP_8970_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3436/do_while_stmt_3437/$exit
      -- 
    timerDaemon_CP_8970_elements(44) <= timerDaemon_CP_8970_elements(3);
    timerDaemon_do_while_stmt_3437_terminator_9085: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_3437_terminator_9085", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_8970_elements(6),loop_continue => timerDaemon_CP_8970_elements(43),loop_terminate => timerDaemon_CP_8970_elements(42),loop_back => timerDaemon_CP_8970_elements(4),loop_exit => timerDaemon_CP_8970_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_3439_phi_seq_9043_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_8970_elements(21);
      timerDaemon_CP_8970_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_8970_elements(24);
      timerDaemon_CP_8970_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_8970_elements(26);
      timerDaemon_CP_8970_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_8970_elements(19);
      timerDaemon_CP_8970_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_8970_elements(30);
      timerDaemon_CP_8970_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_8970_elements(31);
      timerDaemon_CP_8970_elements(20) <= phi_mux_reqs(1);
      phi_stmt_3439_phi_seq_9043 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_3439_phi_seq_9043") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_8970_elements(11), 
          phi_sample_ack => timerDaemon_CP_8970_elements(17), 
          phi_update_req => timerDaemon_CP_8970_elements(13), 
          phi_update_ack => timerDaemon_CP_8970_elements(18), 
          phi_mux_ack => timerDaemon_CP_8970_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_8995_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_8970_elements(7);
        preds(1)  <= timerDaemon_CP_8970_elements(8);
        entry_tmerge_8995 : transition_merge -- 
          generic map(name => " entry_tmerge_8995")
          port map (preds => preds, symbol_out => timerDaemon_CP_8970_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_3439 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_3446_wire : std_logic_vector(0 downto 0);
    signal konst_3450_wire_constant : std_logic_vector(63 downto 0);
    signal konst_3458_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_3452 : std_logic_vector(63 downto 0);
    signal nCOUNTER_3452_3443_buffered : std_logic_vector(63 downto 0);
    signal req_3444 : std_logic_vector(0 downto 0);
    signal type_cast_3442_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_3450_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_3458_wire_constant <= "1";
    type_cast_3442_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_3439: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3442_wire_constant & nCOUNTER_3452_3443_buffered;
      req <= phi_stmt_3439_req_0 & phi_stmt_3439_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3439",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3439_ack_0,
          idata => idata,
          odata => COUNTER_3439,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3439
    nCOUNTER_3452_3443_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_3452_3443_buf_req_0;
      nCOUNTER_3452_3443_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_3452_3443_buf_req_1;
      nCOUNTER_3452_3443_buf_ack_1<= rack(0);
      nCOUNTER_3452_3443_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_3452_3443_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_3452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_3452_3443_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_3444
    process(RPIPE_timer_req_3446_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_3446_wire(0 downto 0);
      req_3444 <= tmp_var; -- 
    end process;
    do_while_stmt_3437_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_3458_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3437_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3437_branch_req_0,
          ack0 => do_while_stmt_3437_branch_ack_0,
          ack1 => do_while_stmt_3437_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_3451_inst
    process(COUNTER_3439) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_3439, konst_3450_wire_constant, tmp_var);
      nCOUNTER_3452 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_3446_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_3446_inst_req_0;
      RPIPE_timer_req_3446_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_3446_inst_req_1;
      RPIPE_timer_req_3446_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_3446_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_3454_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_3454_inst_req_0;
      WPIPE_timer_resp_3454_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_3454_inst_req_1;
      WPIPE_timer_resp_3454_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_3444(0);
      data_in <= COUNTER_3439;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(27 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(27 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(127 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_row_in :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(47 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(47 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(47 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(63 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_num_chl :  std_logic_vector(15 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(79 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(79 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(63 downto 0);
  signal sendB_in_args    : std_logic_vector(63 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(63 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendModule
  component sendModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
      output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendModule
  signal sendModule_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendModule_tag_out   : std_logic_vector(1 downto 0);
  signal sendModule_start_req : std_logic;
  signal sendModule_start_ack : std_logic;
  signal sendModule_fin_req   : std_logic;
  signal sendModule_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe2
  signal input_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe2
  signal input_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe3
  signal input_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe3
  signal input_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe3
  signal kernel_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe3
  signal kernel_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe output_pipe
  signal output_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe output_pipe
  signal output_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_row_in <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 48,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      row_in => access_T_row_in,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(19 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      input_pipe2_pipe_write_req => input_pipe2_pipe_write_req(0 downto 0),
      input_pipe2_pipe_write_ack => input_pipe2_pipe_write_ack(0 downto 0),
      input_pipe2_pipe_write_data => input_pipe2_pipe_write_data(15 downto 0),
      input_pipe3_pipe_write_req => input_pipe3_pipe_write_req(0 downto 0),
      input_pipe3_pipe_write_ack => input_pipe3_pipe_write_ack(0 downto 0),
      input_pipe3_pipe_write_data => input_pipe3_pipe_write_data(15 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(27 downto 14),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(19 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(7 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(1 downto 1),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(1 downto 1),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(31 downto 16),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(47 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(79 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(63 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe2_pipe_read_req => input_pipe2_pipe_read_req(0 downto 0),
      input_pipe2_pipe_read_ack => input_pipe2_pipe_read_ack(0 downto 0),
      input_pipe2_pipe_read_data => input_pipe2_pipe_read_data(15 downto 0),
      input_pipe3_pipe_read_req => input_pipe3_pipe_read_req(0 downto 0),
      input_pipe3_pipe_read_ack => input_pipe3_pipe_read_ack(0 downto 0),
      input_pipe3_pipe_read_data => input_pipe3_pipe_read_data(15 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(15 downto 0),
      kernel_pipe3_pipe_read_req => kernel_pipe3_pipe_read_req(0 downto 0),
      kernel_pipe3_pipe_read_ack => kernel_pipe3_pipe_read_ack(0 downto 0),
      kernel_pipe3_pipe_read_data => kernel_pipe3_pipe_read_data(15 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(1 downto 1),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(1 downto 1),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(15 downto 8),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(0 downto 0),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(0 downto 0),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(79 downto 16);
  loadKernelChannel_num_chl <= loadKernelChannel_in_args(15 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 80,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      num_chl => loadKernelChannel_num_chl,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(1 downto 1),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(1 downto 1),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(15 downto 8),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(15 downto 0),
      kernel_pipe3_pipe_write_req => kernel_pipe3_pipe_write_req(0 downto 0),
      kernel_pipe3_pipe_write_ack => kernel_pipe3_pipe_write_ack(0 downto 0),
      kernel_pipe3_pipe_write_data => kernel_pipe3_pipe_write_data(15 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(15 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(63 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module sendModule
  sendModule_instance:sendModule-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendModule_start_req,
      start_ack => sendModule_start_ack,
      fin_req => sendModule_fin_req,
      fin_ack => sendModule_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      output_pipe_pipe_read_req => output_pipe_pipe_read_req(1 downto 0),
      output_pipe_pipe_read_ack => output_pipe_pipe_read_ack(1 downto 0),
      output_pipe_pipe_read_data => output_pipe_pipe_read_data(31 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(7 downto 0),
      tag_in => sendModule_tag_in,
      tag_out => sendModule_tag_out-- 
    ); -- 
  -- module will be run forever 
  sendModule_tag_in <= (others => '0');
  sendModule_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => sendModule_start_req, start_ack => sendModule_start_ack,  fin_req => sendModule_fin_req,  fin_ack => sendModule_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe2_pipe_read_req,
      read_ack => input_pipe2_pipe_read_ack,
      read_data => input_pipe2_pipe_read_data,
      write_req => input_pipe2_pipe_write_req,
      write_ack => input_pipe2_pipe_write_ack,
      write_data => input_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe3_pipe_read_req,
      read_ack => input_pipe3_pipe_read_ack,
      read_data => input_pipe3_pipe_read_data,
      write_req => input_pipe3_pipe_write_req,
      write_ack => input_pipe3_pipe_write_ack,
      write_data => input_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe3_pipe_read_req,
      read_ack => kernel_pipe3_pipe_read_ack,
      read_data => kernel_pipe3_pipe_read_data,
      write_req => kernel_pipe3_pipe_write_req,
      write_ack => kernel_pipe3_pipe_write_ack,
      write_data => kernel_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe output_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 10 --
    )
    port map( -- 
      read_req => output_pipe_pipe_read_req,
      read_ack => output_pipe_pipe_read_ack,
      read_data => output_pipe_pipe_read_data,
      write_req => output_pipe_pipe_write_req,
      write_ack => output_pipe_pipe_write_ack,
      write_data => output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 11 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 2,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
