-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity concat is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
    Concat_input_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
    Concat_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity concat;
architecture concat_arch of concat is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal concat_CP_34_start: Boolean;
  signal concat_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_Concat_input_pipe_619_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_655_inst_ack_1 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_ack_0 : boolean;
  signal type_cast_641_inst_req_0 : boolean;
  signal type_cast_473_inst_ack_1 : boolean;
  signal if_stmt_537_branch_ack_1 : boolean;
  signal addr_of_603_final_reg_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_ack_0 : boolean;
  signal type_cast_473_inst_req_1 : boolean;
  signal type_cast_509_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_487_inst_ack_1 : boolean;
  signal type_cast_473_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_487_inst_req_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_ack_1 : boolean;
  signal type_cast_1270_inst_req_0 : boolean;
  signal type_cast_837_inst_req_1 : boolean;
  signal type_cast_30_inst_req_0 : boolean;
  signal type_cast_30_inst_ack_0 : boolean;
  signal type_cast_30_inst_req_1 : boolean;
  signal type_cast_30_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_655_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_ack_1 : boolean;
  signal phi_stmt_839_req_0 : boolean;
  signal type_cast_43_inst_req_0 : boolean;
  signal type_cast_43_inst_ack_0 : boolean;
  signal type_cast_43_inst_req_1 : boolean;
  signal type_cast_43_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_655_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_ack_0 : boolean;
  signal type_cast_610_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_606_inst_ack_0 : boolean;
  signal phi_stmt_839_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_req_1 : boolean;
  signal if_stmt_537_branch_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_606_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_637_inst_req_0 : boolean;
  signal type_cast_847_inst_ack_0 : boolean;
  signal type_cast_55_inst_req_0 : boolean;
  signal type_cast_55_inst_ack_0 : boolean;
  signal type_cast_847_inst_req_1 : boolean;
  signal type_cast_55_inst_req_1 : boolean;
  signal type_cast_55_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_ack_0 : boolean;
  signal type_cast_509_inst_req_1 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_ack_1 : boolean;
  signal type_cast_68_inst_req_0 : boolean;
  signal type_cast_68_inst_ack_0 : boolean;
  signal type_cast_68_inst_req_1 : boolean;
  signal type_cast_68_inst_ack_1 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_606_inst_req_1 : boolean;
  signal type_cast_80_inst_req_0 : boolean;
  signal type_cast_80_inst_ack_0 : boolean;
  signal type_cast_595_inst_ack_1 : boolean;
  signal type_cast_80_inst_req_1 : boolean;
  signal type_cast_80_inst_ack_1 : boolean;
  signal type_cast_847_inst_req_0 : boolean;
  signal type_cast_509_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_ack_1 : boolean;
  signal type_cast_1171_inst_req_1 : boolean;
  signal type_cast_93_inst_req_0 : boolean;
  signal type_cast_93_inst_ack_0 : boolean;
  signal type_cast_595_inst_req_1 : boolean;
  signal type_cast_93_inst_req_1 : boolean;
  signal type_cast_93_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_ack_0 : boolean;
  signal type_cast_509_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_ack_1 : boolean;
  signal type_cast_105_inst_req_0 : boolean;
  signal type_cast_105_inst_ack_0 : boolean;
  signal type_cast_105_inst_req_1 : boolean;
  signal type_cast_105_inst_ack_1 : boolean;
  signal array_obj_ref_602_index_offset_ack_1 : boolean;
  signal array_obj_ref_602_index_offset_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_ack_1 : boolean;
  signal type_cast_118_inst_req_0 : boolean;
  signal type_cast_1171_inst_ack_0 : boolean;
  signal type_cast_118_inst_ack_0 : boolean;
  signal type_cast_595_inst_ack_0 : boolean;
  signal type_cast_118_inst_req_1 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_req_1 : boolean;
  signal type_cast_118_inst_ack_1 : boolean;
  signal ptr_deref_1543_load_0_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_req_0 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_ack_1 : boolean;
  signal type_cast_130_inst_req_0 : boolean;
  signal type_cast_130_inst_ack_0 : boolean;
  signal type_cast_595_inst_req_0 : boolean;
  signal type_cast_130_inst_req_1 : boolean;
  signal type_cast_130_inst_ack_1 : boolean;
  signal type_cast_837_inst_ack_0 : boolean;
  signal array_obj_ref_602_index_offset_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_619_inst_ack_0 : boolean;
  signal MUX_1253_inst_ack_1 : boolean;
  signal ptr_deref_517_store_0_ack_0 : boolean;
  signal ptr_deref_517_store_0_req_0 : boolean;
  signal ptr_deref_885_load_0_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_619_inst_req_1 : boolean;
  signal type_cast_143_inst_req_0 : boolean;
  signal type_cast_143_inst_ack_0 : boolean;
  signal type_cast_143_inst_req_1 : boolean;
  signal type_cast_143_inst_ack_1 : boolean;
  signal array_obj_ref_602_index_offset_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_ack_0 : boolean;
  signal type_cast_610_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_req_1 : boolean;
  signal do_while_stmt_368_branch_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_ack_1 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal ptr_deref_885_load_0_req_1 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_606_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_637_inst_ack_0 : boolean;
  signal type_cast_837_inst_ack_1 : boolean;
  signal type_cast_168_inst_req_0 : boolean;
  signal do_while_stmt_368_branch_ack_0 : boolean;
  signal type_cast_168_inst_ack_0 : boolean;
  signal type_cast_168_inst_req_1 : boolean;
  signal type_cast_168_inst_ack_1 : boolean;
  signal type_cast_837_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_ack_0 : boolean;
  signal type_cast_610_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_ack_1 : boolean;
  signal type_cast_567_inst_ack_1 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_0 : boolean;
  signal type_cast_180_inst_req_0 : boolean;
  signal type_cast_180_inst_ack_0 : boolean;
  signal ptr_deref_885_load_0_ack_1 : boolean;
  signal type_cast_180_inst_req_1 : boolean;
  signal type_cast_1171_inst_req_0 : boolean;
  signal type_cast_180_inst_ack_1 : boolean;
  signal type_cast_623_inst_ack_1 : boolean;
  signal type_cast_567_inst_req_1 : boolean;
  signal type_cast_610_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_505_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_ack_1 : boolean;
  signal type_cast_193_inst_req_0 : boolean;
  signal type_cast_193_inst_ack_0 : boolean;
  signal type_cast_193_inst_req_1 : boolean;
  signal type_cast_193_inst_ack_1 : boolean;
  signal type_cast_623_inst_req_1 : boolean;
  signal phi_stmt_839_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_505_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_637_inst_ack_1 : boolean;
  signal type_cast_567_inst_ack_0 : boolean;
  signal type_cast_205_inst_req_0 : boolean;
  signal type_cast_205_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_req_1 : boolean;
  signal type_cast_205_inst_req_1 : boolean;
  signal type_cast_205_inst_ack_1 : boolean;
  signal type_cast_641_inst_ack_1 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_637_inst_req_1 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_req_1 : boolean;
  signal type_cast_567_inst_req_0 : boolean;
  signal ptr_deref_517_store_0_ack_1 : boolean;
  signal type_cast_218_inst_req_0 : boolean;
  signal type_cast_473_inst_req_0 : boolean;
  signal type_cast_218_inst_ack_0 : boolean;
  signal type_cast_218_inst_req_1 : boolean;
  signal type_cast_218_inst_ack_1 : boolean;
  signal type_cast_641_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_ack_1 : boolean;
  signal ptr_deref_517_store_0_req_1 : boolean;
  signal type_cast_230_inst_req_0 : boolean;
  signal type_cast_230_inst_ack_0 : boolean;
  signal type_cast_230_inst_req_1 : boolean;
  signal type_cast_230_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_505_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_ack_1 : boolean;
  signal type_cast_243_inst_req_0 : boolean;
  signal type_cast_243_inst_ack_0 : boolean;
  signal type_cast_243_inst_req_1 : boolean;
  signal type_cast_243_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_505_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_487_inst_ack_0 : boolean;
  signal if_stmt_298_branch_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_487_inst_req_0 : boolean;
  signal if_stmt_298_branch_ack_1 : boolean;
  signal if_stmt_298_branch_ack_0 : boolean;
  signal if_stmt_313_branch_req_0 : boolean;
  signal if_stmt_313_branch_ack_1 : boolean;
  signal if_stmt_313_branch_ack_0 : boolean;
  signal array_obj_ref_899_index_offset_req_0 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal type_cast_623_inst_ack_0 : boolean;
  signal type_cast_641_inst_ack_0 : boolean;
  signal do_while_stmt_368_branch_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_619_inst_ack_1 : boolean;
  signal type_cast_1186_inst_req_0 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_ack_1 : boolean;
  signal phi_stmt_592_ack_0 : boolean;
  signal addr_of_603_final_reg_ack_1 : boolean;
  signal phi_stmt_370_req_0 : boolean;
  signal type_cast_847_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_655_inst_req_1 : boolean;
  signal phi_stmt_370_req_1 : boolean;
  signal phi_stmt_370_ack_0 : boolean;
  signal addr_of_603_final_reg_req_1 : boolean;
  signal type_cast_373_inst_req_0 : boolean;
  signal type_cast_373_inst_ack_0 : boolean;
  signal type_cast_373_inst_req_1 : boolean;
  signal type_cast_373_inst_ack_1 : boolean;
  signal type_cast_623_inst_req_0 : boolean;
  signal phi_stmt_592_req_0 : boolean;
  signal do_while_stmt_590_branch_req_0 : boolean;
  signal array_obj_ref_380_index_offset_req_0 : boolean;
  signal array_obj_ref_380_index_offset_ack_0 : boolean;
  signal array_obj_ref_380_index_offset_req_1 : boolean;
  signal array_obj_ref_380_index_offset_ack_1 : boolean;
  signal type_cast_491_inst_ack_1 : boolean;
  signal type_cast_491_inst_req_1 : boolean;
  signal phi_stmt_592_req_1 : boolean;
  signal addr_of_381_final_reg_req_0 : boolean;
  signal addr_of_381_final_reg_ack_0 : boolean;
  signal addr_of_381_final_reg_req_1 : boolean;
  signal addr_of_381_final_reg_ack_1 : boolean;
  signal type_cast_491_inst_ack_0 : boolean;
  signal addr_of_603_final_reg_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_384_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_384_inst_ack_0 : boolean;
  signal type_cast_491_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_384_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_384_inst_ack_1 : boolean;
  signal type_cast_388_inst_req_0 : boolean;
  signal type_cast_388_inst_ack_0 : boolean;
  signal type_cast_388_inst_req_1 : boolean;
  signal type_cast_388_inst_ack_1 : boolean;
  signal if_stmt_537_branch_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_397_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_397_inst_ack_0 : boolean;
  signal type_cast_870_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_397_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_397_inst_ack_1 : boolean;
  signal type_cast_870_inst_ack_0 : boolean;
  signal MUX_1253_inst_req_0 : boolean;
  signal type_cast_401_inst_req_0 : boolean;
  signal type_cast_401_inst_ack_0 : boolean;
  signal type_cast_401_inst_req_1 : boolean;
  signal type_cast_401_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_req_0 : boolean;
  signal ptr_deref_885_load_0_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_415_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_415_inst_ack_0 : boolean;
  signal type_cast_870_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_415_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_415_inst_ack_1 : boolean;
  signal type_cast_870_inst_ack_1 : boolean;
  signal type_cast_419_inst_req_0 : boolean;
  signal type_cast_419_inst_ack_0 : boolean;
  signal type_cast_419_inst_req_1 : boolean;
  signal type_cast_419_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_433_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_433_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_433_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_433_inst_ack_1 : boolean;
  signal type_cast_437_inst_req_0 : boolean;
  signal type_cast_437_inst_ack_0 : boolean;
  signal type_cast_437_inst_req_1 : boolean;
  signal type_cast_437_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_451_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_451_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_451_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_451_inst_ack_1 : boolean;
  signal type_cast_455_inst_req_0 : boolean;
  signal type_cast_455_inst_ack_0 : boolean;
  signal type_cast_455_inst_req_1 : boolean;
  signal type_cast_455_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_469_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_469_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_469_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_469_inst_ack_1 : boolean;
  signal type_cast_659_inst_req_0 : boolean;
  signal type_cast_659_inst_ack_0 : boolean;
  signal type_cast_659_inst_req_1 : boolean;
  signal type_cast_659_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_673_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_673_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_673_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_673_inst_ack_1 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_1 : boolean;
  signal type_cast_893_inst_ack_1 : boolean;
  signal type_cast_677_inst_req_0 : boolean;
  signal type_cast_677_inst_ack_0 : boolean;
  signal type_cast_677_inst_req_1 : boolean;
  signal type_cast_677_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_ack_0 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_691_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_691_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_691_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_691_inst_ack_1 : boolean;
  signal type_cast_695_inst_req_0 : boolean;
  signal type_cast_695_inst_ack_0 : boolean;
  signal type_cast_695_inst_req_1 : boolean;
  signal type_cast_695_inst_ack_1 : boolean;
  signal MUX_1253_inst_ack_0 : boolean;
  signal W_arrayidx245_894_delayed_6_0_905_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_709_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_709_inst_ack_0 : boolean;
  signal W_arrayidx245_894_delayed_6_0_905_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_709_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_709_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_0 : boolean;
  signal type_cast_893_inst_req_1 : boolean;
  signal type_cast_1270_inst_ack_0 : boolean;
  signal array_obj_ref_899_index_offset_ack_1 : boolean;
  signal type_cast_713_inst_req_0 : boolean;
  signal type_cast_1171_inst_ack_1 : boolean;
  signal type_cast_713_inst_ack_0 : boolean;
  signal type_cast_713_inst_req_1 : boolean;
  signal type_cast_713_inst_ack_1 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_0 : boolean;
  signal ptr_deref_910_store_0_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_727_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_727_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_727_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_727_inst_ack_1 : boolean;
  signal array_obj_ref_899_index_offset_req_1 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_1 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal type_cast_731_inst_req_0 : boolean;
  signal type_cast_731_inst_ack_0 : boolean;
  signal type_cast_731_inst_req_1 : boolean;
  signal type_cast_731_inst_ack_1 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_0 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_0 : boolean;
  signal type_cast_842_inst_ack_1 : boolean;
  signal addr_of_877_final_reg_ack_1 : boolean;
  signal addr_of_877_final_reg_req_1 : boolean;
  signal type_cast_1270_inst_ack_1 : boolean;
  signal W_arrayidx245_894_delayed_6_0_905_inst_ack_0 : boolean;
  signal ptr_deref_739_store_0_req_0 : boolean;
  signal ptr_deref_739_store_0_ack_0 : boolean;
  signal ptr_deref_739_store_0_req_1 : boolean;
  signal addr_of_877_final_reg_ack_0 : boolean;
  signal ptr_deref_739_store_0_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_ack_1 : boolean;
  signal addr_of_877_final_reg_req_0 : boolean;
  signal type_cast_842_inst_req_1 : boolean;
  signal type_cast_893_inst_ack_0 : boolean;
  signal W_arrayidx245_894_delayed_6_0_905_inst_req_0 : boolean;
  signal array_obj_ref_876_index_offset_ack_1 : boolean;
  signal array_obj_ref_876_index_offset_req_1 : boolean;
  signal addr_of_900_final_reg_ack_1 : boolean;
  signal type_cast_893_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_req_1 : boolean;
  signal do_while_stmt_590_branch_ack_0 : boolean;
  signal do_while_stmt_590_branch_ack_1 : boolean;
  signal array_obj_ref_876_index_offset_ack_0 : boolean;
  signal ptr_deref_910_store_0_ack_0 : boolean;
  signal type_cast_842_inst_ack_0 : boolean;
  signal array_obj_ref_899_index_offset_ack_0 : boolean;
  signal if_stmt_759_branch_req_0 : boolean;
  signal if_stmt_759_branch_ack_1 : boolean;
  signal if_stmt_759_branch_ack_0 : boolean;
  signal type_cast_842_inst_req_0 : boolean;
  signal array_obj_ref_876_index_offset_req_0 : boolean;
  signal call_stmt_768_call_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_req_1 : boolean;
  signal call_stmt_768_call_ack_0 : boolean;
  signal call_stmt_768_call_req_1 : boolean;
  signal call_stmt_768_call_ack_1 : boolean;
  signal addr_of_900_final_reg_req_1 : boolean;
  signal do_while_stmt_817_branch_req_0 : boolean;
  signal MUX_1253_inst_req_1 : boolean;
  signal addr_of_900_final_reg_ack_0 : boolean;
  signal type_cast_1274_inst_req_0 : boolean;
  signal phi_stmt_819_req_0 : boolean;
  signal addr_of_900_final_reg_req_0 : boolean;
  signal phi_stmt_819_req_1 : boolean;
  signal type_cast_1242_inst_req_0 : boolean;
  signal phi_stmt_819_ack_0 : boolean;
  signal type_cast_1242_inst_ack_0 : boolean;
  signal type_cast_1186_inst_ack_0 : boolean;
  signal type_cast_1242_inst_req_1 : boolean;
  signal type_cast_1202_inst_req_0 : boolean;
  signal type_cast_822_inst_req_0 : boolean;
  signal type_cast_822_inst_ack_0 : boolean;
  signal type_cast_1202_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_1 : boolean;
  signal type_cast_822_inst_ack_1 : boolean;
  signal type_cast_1242_inst_ack_1 : boolean;
  signal type_cast_1266_inst_req_1 : boolean;
  signal type_cast_1274_inst_req_1 : boolean;
  signal type_cast_1274_inst_ack_0 : boolean;
  signal phi_stmt_824_req_0 : boolean;
  signal type_cast_1274_inst_ack_1 : boolean;
  signal phi_stmt_824_req_1 : boolean;
  signal type_cast_1270_inst_req_1 : boolean;
  signal phi_stmt_824_ack_0 : boolean;
  signal type_cast_1246_inst_req_0 : boolean;
  signal type_cast_1246_inst_ack_0 : boolean;
  signal type_cast_827_inst_req_0 : boolean;
  signal type_cast_827_inst_ack_0 : boolean;
  signal type_cast_827_inst_req_1 : boolean;
  signal type_cast_827_inst_ack_1 : boolean;
  signal type_cast_1186_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_ack_0 : boolean;
  signal type_cast_1246_inst_req_1 : boolean;
  signal type_cast_1246_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_ack_0 : boolean;
  signal type_cast_1266_inst_ack_1 : boolean;
  signal array_obj_ref_1538_index_offset_req_0 : boolean;
  signal phi_stmt_829_req_0 : boolean;
  signal phi_stmt_829_req_1 : boolean;
  signal phi_stmt_829_ack_0 : boolean;
  signal type_cast_832_inst_req_0 : boolean;
  signal type_cast_832_inst_ack_0 : boolean;
  signal type_cast_832_inst_req_1 : boolean;
  signal type_cast_832_inst_ack_1 : boolean;
  signal phi_stmt_834_req_0 : boolean;
  signal phi_stmt_834_req_1 : boolean;
  signal phi_stmt_834_ack_0 : boolean;
  signal array_obj_ref_1538_index_offset_ack_0 : boolean;
  signal type_cast_1266_inst_req_0 : boolean;
  signal type_cast_1266_inst_ack_0 : boolean;
  signal ptr_deref_910_store_0_req_1 : boolean;
  signal W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_req_0 : boolean;
  signal ptr_deref_910_store_0_ack_1 : boolean;
  signal type_cast_1202_inst_ack_1 : boolean;
  signal type_cast_1202_inst_req_1 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_req_0 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_0 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_req_1 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_req_0 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_req_0 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_0 : boolean;
  signal type_cast_1186_inst_ack_1 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_req_1 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_ack_0 : boolean;
  signal type_cast_1509_inst_req_0 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_req_0 : boolean;
  signal type_cast_1509_inst_ack_0 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_ack_0 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_req_1 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_req_1 : boolean;
  signal type_cast_1587_inst_req_0 : boolean;
  signal type_cast_953_inst_req_0 : boolean;
  signal type_cast_953_inst_ack_0 : boolean;
  signal type_cast_1587_inst_ack_0 : boolean;
  signal type_cast_953_inst_req_1 : boolean;
  signal type_cast_953_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_ack_1 : boolean;
  signal type_cast_968_inst_req_0 : boolean;
  signal type_cast_968_inst_ack_0 : boolean;
  signal type_cast_968_inst_req_1 : boolean;
  signal type_cast_968_inst_ack_1 : boolean;
  signal type_cast_1509_inst_req_1 : boolean;
  signal type_cast_1567_inst_req_0 : boolean;
  signal type_cast_1509_inst_ack_1 : boolean;
  signal type_cast_983_inst_req_0 : boolean;
  signal type_cast_983_inst_ack_0 : boolean;
  signal type_cast_983_inst_req_1 : boolean;
  signal type_cast_983_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_req_1 : boolean;
  signal type_cast_1567_inst_ack_0 : boolean;
  signal type_cast_1597_inst_ack_1 : boolean;
  signal type_cast_1597_inst_req_1 : boolean;
  signal type_cast_999_inst_req_0 : boolean;
  signal type_cast_999_inst_ack_0 : boolean;
  signal array_obj_ref_1538_index_offset_req_1 : boolean;
  signal type_cast_1587_inst_req_1 : boolean;
  signal type_cast_999_inst_req_1 : boolean;
  signal type_cast_999_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_req_0 : boolean;
  signal array_obj_ref_1538_index_offset_ack_1 : boolean;
  signal type_cast_1567_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_1 : boolean;
  signal type_cast_1587_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_ack_0 : boolean;
  signal type_cast_1567_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_1 : boolean;
  signal type_cast_1547_inst_req_0 : boolean;
  signal type_cast_1547_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_1 : boolean;
  signal type_cast_1547_inst_req_1 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_0 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_0 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_1 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_req_0 : boolean;
  signal type_cast_1036_inst_req_0 : boolean;
  signal type_cast_1036_inst_ack_0 : boolean;
  signal type_cast_1036_inst_req_1 : boolean;
  signal type_cast_1036_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_ack_0 : boolean;
  signal type_cast_1547_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_req_0 : boolean;
  signal type_cast_1577_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_req_1 : boolean;
  signal type_cast_1577_inst_ack_0 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_0 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_0 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_1 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_ack_0 : boolean;
  signal type_cast_1597_inst_req_0 : boolean;
  signal ptr_deref_1543_load_0_req_0 : boolean;
  signal type_cast_1557_inst_req_0 : boolean;
  signal type_cast_1073_inst_req_0 : boolean;
  signal type_cast_1073_inst_ack_0 : boolean;
  signal type_cast_1073_inst_req_1 : boolean;
  signal type_cast_1073_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_ack_1 : boolean;
  signal type_cast_1557_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_req_1 : boolean;
  signal ptr_deref_1543_load_0_ack_0 : boolean;
  signal array_obj_ref_1079_index_offset_req_0 : boolean;
  signal array_obj_ref_1079_index_offset_ack_0 : boolean;
  signal array_obj_ref_1079_index_offset_req_1 : boolean;
  signal array_obj_ref_1079_index_offset_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_ack_0 : boolean;
  signal addr_of_1080_final_reg_req_0 : boolean;
  signal addr_of_1080_final_reg_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_ack_1 : boolean;
  signal addr_of_1080_final_reg_req_1 : boolean;
  signal addr_of_1080_final_reg_ack_1 : boolean;
  signal W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_req_0 : boolean;
  signal W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_ack_0 : boolean;
  signal W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_req_1 : boolean;
  signal W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_ack_1 : boolean;
  signal ptr_deref_1088_load_0_req_0 : boolean;
  signal ptr_deref_1088_load_0_ack_0 : boolean;
  signal ptr_deref_1088_load_0_req_1 : boolean;
  signal ptr_deref_1088_load_0_ack_1 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_req_0 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_0 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_req_1 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_1 : boolean;
  signal type_cast_1096_inst_req_0 : boolean;
  signal type_cast_1096_inst_ack_0 : boolean;
  signal type_cast_1096_inst_req_1 : boolean;
  signal type_cast_1096_inst_ack_1 : boolean;
  signal array_obj_ref_1102_index_offset_req_0 : boolean;
  signal array_obj_ref_1102_index_offset_ack_0 : boolean;
  signal array_obj_ref_1102_index_offset_req_1 : boolean;
  signal array_obj_ref_1102_index_offset_ack_1 : boolean;
  signal addr_of_1103_final_reg_req_0 : boolean;
  signal addr_of_1103_final_reg_ack_0 : boolean;
  signal addr_of_1103_final_reg_req_1 : boolean;
  signal addr_of_1103_final_reg_ack_1 : boolean;
  signal W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_req_0 : boolean;
  signal W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_ack_0 : boolean;
  signal W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_req_1 : boolean;
  signal W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_ack_1 : boolean;
  signal W_arrayidx273_1043_delayed_6_0_1108_inst_req_0 : boolean;
  signal W_arrayidx273_1043_delayed_6_0_1108_inst_ack_0 : boolean;
  signal W_arrayidx273_1043_delayed_6_0_1108_inst_req_1 : boolean;
  signal W_arrayidx273_1043_delayed_6_0_1108_inst_ack_1 : boolean;
  signal ptr_deref_1113_store_0_req_0 : boolean;
  signal ptr_deref_1113_store_0_ack_0 : boolean;
  signal ptr_deref_1113_store_0_req_1 : boolean;
  signal ptr_deref_1113_store_0_ack_1 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_0 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_0 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_1 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_1 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_0 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_0 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_1 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_1 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_req_0 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_0 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_req_1 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_1 : boolean;
  signal type_cast_1156_inst_req_0 : boolean;
  signal type_cast_1156_inst_ack_0 : boolean;
  signal type_cast_1156_inst_req_1 : boolean;
  signal type_cast_1156_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_req_0 : boolean;
  signal MUX_1281_inst_req_0 : boolean;
  signal MUX_1281_inst_ack_0 : boolean;
  signal MUX_1281_inst_req_1 : boolean;
  signal MUX_1281_inst_ack_1 : boolean;
  signal ptr_deref_1543_load_0_req_1 : boolean;
  signal type_cast_1597_inst_ack_0 : boolean;
  signal type_cast_1557_inst_ack_1 : boolean;
  signal type_cast_1557_inst_req_1 : boolean;
  signal if_stmt_1488_branch_ack_0 : boolean;
  signal addr_of_1539_final_reg_ack_1 : boolean;
  signal if_stmt_1488_branch_ack_1 : boolean;
  signal type_cast_1294_inst_req_0 : boolean;
  signal addr_of_1539_final_reg_req_1 : boolean;
  signal type_cast_1294_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_ack_1 : boolean;
  signal type_cast_1294_inst_req_1 : boolean;
  signal type_cast_1294_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_req_1 : boolean;
  signal if_stmt_1488_branch_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_req_1 : boolean;
  signal type_cast_1577_inst_ack_1 : boolean;
  signal type_cast_1298_inst_req_0 : boolean;
  signal addr_of_1539_final_reg_ack_0 : boolean;
  signal type_cast_1298_inst_ack_0 : boolean;
  signal type_cast_1577_inst_req_1 : boolean;
  signal type_cast_1298_inst_req_1 : boolean;
  signal addr_of_1539_final_reg_req_0 : boolean;
  signal type_cast_1298_inst_ack_1 : boolean;
  signal MUX_1305_inst_req_0 : boolean;
  signal MUX_1305_inst_ack_0 : boolean;
  signal MUX_1305_inst_req_1 : boolean;
  signal MUX_1305_inst_ack_1 : boolean;
  signal type_cast_1320_inst_req_0 : boolean;
  signal type_cast_1320_inst_ack_0 : boolean;
  signal type_cast_1320_inst_req_1 : boolean;
  signal type_cast_1320_inst_ack_1 : boolean;
  signal type_cast_1324_inst_req_0 : boolean;
  signal type_cast_1324_inst_ack_0 : boolean;
  signal type_cast_1324_inst_req_1 : boolean;
  signal type_cast_1324_inst_ack_1 : boolean;
  signal MUX_1331_inst_req_0 : boolean;
  signal MUX_1331_inst_ack_0 : boolean;
  signal MUX_1331_inst_req_1 : boolean;
  signal MUX_1331_inst_ack_1 : boolean;
  signal type_cast_1346_inst_req_0 : boolean;
  signal type_cast_1346_inst_ack_0 : boolean;
  signal type_cast_1346_inst_req_1 : boolean;
  signal type_cast_1346_inst_ack_1 : boolean;
  signal do_while_stmt_817_branch_ack_0 : boolean;
  signal do_while_stmt_817_branch_ack_1 : boolean;
  signal if_stmt_1359_branch_req_0 : boolean;
  signal if_stmt_1359_branch_ack_1 : boolean;
  signal if_stmt_1359_branch_ack_0 : boolean;
  signal type_cast_1368_inst_req_0 : boolean;
  signal type_cast_1368_inst_ack_0 : boolean;
  signal type_cast_1368_inst_req_1 : boolean;
  signal type_cast_1368_inst_ack_1 : boolean;
  signal call_stmt_1372_call_req_0 : boolean;
  signal call_stmt_1372_call_ack_0 : boolean;
  signal call_stmt_1372_call_req_1 : boolean;
  signal call_stmt_1372_call_ack_1 : boolean;
  signal type_cast_1376_inst_req_0 : boolean;
  signal type_cast_1376_inst_ack_0 : boolean;
  signal type_cast_1376_inst_req_1 : boolean;
  signal type_cast_1376_inst_ack_1 : boolean;
  signal type_cast_1385_inst_req_0 : boolean;
  signal type_cast_1385_inst_ack_0 : boolean;
  signal type_cast_1385_inst_req_1 : boolean;
  signal type_cast_1385_inst_ack_1 : boolean;
  signal type_cast_1395_inst_req_0 : boolean;
  signal type_cast_1395_inst_ack_0 : boolean;
  signal type_cast_1395_inst_req_1 : boolean;
  signal type_cast_1395_inst_ack_1 : boolean;
  signal type_cast_1405_inst_req_0 : boolean;
  signal type_cast_1405_inst_ack_0 : boolean;
  signal type_cast_1405_inst_req_1 : boolean;
  signal type_cast_1405_inst_ack_1 : boolean;
  signal type_cast_1415_inst_req_0 : boolean;
  signal type_cast_1415_inst_ack_0 : boolean;
  signal type_cast_1415_inst_req_1 : boolean;
  signal type_cast_1415_inst_ack_1 : boolean;
  signal type_cast_1425_inst_req_0 : boolean;
  signal type_cast_1425_inst_ack_0 : boolean;
  signal type_cast_1425_inst_req_1 : boolean;
  signal type_cast_1425_inst_ack_1 : boolean;
  signal type_cast_1435_inst_req_0 : boolean;
  signal type_cast_1435_inst_ack_0 : boolean;
  signal type_cast_1435_inst_req_1 : boolean;
  signal type_cast_1435_inst_ack_1 : boolean;
  signal type_cast_1445_inst_req_0 : boolean;
  signal type_cast_1445_inst_ack_0 : boolean;
  signal type_cast_1445_inst_req_1 : boolean;
  signal type_cast_1445_inst_ack_1 : boolean;
  signal type_cast_1455_inst_req_0 : boolean;
  signal type_cast_1455_inst_ack_0 : boolean;
  signal type_cast_1455_inst_req_1 : boolean;
  signal type_cast_1455_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_ack_0 : boolean;
  signal type_cast_1607_inst_req_0 : boolean;
  signal type_cast_1607_inst_ack_0 : boolean;
  signal type_cast_1607_inst_req_1 : boolean;
  signal type_cast_1607_inst_ack_1 : boolean;
  signal type_cast_1617_inst_req_0 : boolean;
  signal type_cast_1617_inst_ack_0 : boolean;
  signal type_cast_1617_inst_req_1 : boolean;
  signal type_cast_1617_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_ack_1 : boolean;
  signal if_stmt_1654_branch_req_0 : boolean;
  signal if_stmt_1654_branch_ack_1 : boolean;
  signal if_stmt_1654_branch_ack_0 : boolean;
  signal phi_stmt_1526_req_0 : boolean;
  signal type_cast_1532_inst_req_0 : boolean;
  signal type_cast_1532_inst_ack_0 : boolean;
  signal type_cast_1532_inst_req_1 : boolean;
  signal type_cast_1532_inst_ack_1 : boolean;
  signal phi_stmt_1526_req_1 : boolean;
  signal phi_stmt_1526_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "concat_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  concat_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "concat_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= concat_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  concat_CP_34: Block -- control-path 
    signal concat_CP_34_elements: BooleanArray(802 downto 0);
    -- 
  begin -- 
    concat_CP_34_elements(0) <= concat_CP_34_start;
    concat_CP_34_symbol <= concat_CP_34_elements(802);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	63 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	51 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	43 
    -- CP-element group 0: 	35 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	75 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	31 
    -- CP-element group 0:  members (62) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_23/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/branch_block_stmt_23__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Update/cr
      -- 
    rr_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => RPIPE_Concat_input_pipe_25_inst_req_0); -- 
    cr_143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_30_inst_req_1); -- 
    cr_171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_43_inst_req_1); -- 
    cr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_55_inst_req_1); -- 
    cr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_68_inst_req_1); -- 
    cr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_80_inst_req_1); -- 
    cr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_93_inst_req_1); -- 
    cr_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_105_inst_req_1); -- 
    cr_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_118_inst_req_1); -- 
    cr_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_130_inst_req_1); -- 
    cr_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_143_inst_req_1); -- 
    cr_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_155_inst_req_1); -- 
    cr_451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_168_inst_req_1); -- 
    cr_479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_180_inst_req_1); -- 
    cr_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_193_inst_req_1); -- 
    cr_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_205_inst_req_1); -- 
    cr_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_218_inst_req_1); -- 
    cr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_230_inst_req_1); -- 
    cr_619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_243_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	191 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	192 
    -- CP-element group 1: 	193 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_537_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/do_while_stmt_368__exit__
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_537__entry__
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_537_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/R_forx_xbody_forx_xcond163x_xpreheaderx_xloopexit_taken_538_place
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_537_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_537_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_537_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_537_dead_link/$entry
      -- 
    branch_req_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => if_stmt_537_branch_req_0); -- 
    concat_CP_34_elements(1) <= concat_CP_34_elements(191);
    -- CP-element group 2:  branch  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	304 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	305 
    -- CP-element group 2: 	306 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_23/do_while_stmt_590__exit__
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_759__entry__
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_759_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_759_eval_test/$entry
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_759_eval_test/$exit
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_759_eval_test/branch_req
      -- CP-element group 2: 	 branch_block_stmt_23/R_forx_xbody169_forx_xend223x_xloopexit_taken_760_place
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_759_if_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_759_else_link/$entry
      -- 
    branch_req_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(2), ack => if_stmt_759_branch_req_0); -- 
    concat_CP_34_elements(2) <= concat_CP_34_elements(304);
    -- CP-element group 3:  branch  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	694 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	695 
    -- CP-element group 3: 	696 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_23/do_while_stmt_817__exit__
      -- CP-element group 3: 	 branch_block_stmt_23/if_stmt_1359__entry__
      -- CP-element group 3: 	 branch_block_stmt_23/if_stmt_1359_dead_link/$entry
      -- CP-element group 3: 	 branch_block_stmt_23/if_stmt_1359_eval_test/$entry
      -- CP-element group 3: 	 branch_block_stmt_23/if_stmt_1359_eval_test/$exit
      -- CP-element group 3: 	 branch_block_stmt_23/if_stmt_1359_eval_test/branch_req
      -- CP-element group 3: 	 branch_block_stmt_23/R_ifx_xend297_whilex_xend_taken_1360_place
      -- CP-element group 3: 	 branch_block_stmt_23/if_stmt_1359_if_link/$entry
      -- CP-element group 3: 	 branch_block_stmt_23/if_stmt_1359_else_link/$entry
      -- 
    branch_req_2953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(3), ack => if_stmt_1359_branch_req_0); -- 
    concat_CP_34_elements(3) <= concat_CP_34_elements(694);
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_update_start_
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Update/cr
      -- 
    ra_125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_25_inst_ack_0, ack => concat_CP_34_elements(4)); -- 
    cr_129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(4), ack => RPIPE_Concat_input_pipe_25_inst_req_1); -- 
    -- CP-element group 5:  fork  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_25_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Sample/rr
      -- 
    ca_130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_25_inst_ack_1, ack => concat_CP_34_elements(5)); -- 
    rr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(5), ack => type_cast_30_inst_req_0); -- 
    rr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(5), ack => RPIPE_Concat_input_pipe_39_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Sample/ra
      -- 
    ra_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_30_inst_ack_0, ack => concat_CP_34_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	76 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_30_Update/ca
      -- 
    ca_144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_30_inst_ack_1, ack => concat_CP_34_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_update_start_
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Update/cr
      -- 
    ra_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_39_inst_ack_0, ack => concat_CP_34_elements(8)); -- 
    cr_157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(8), ack => RPIPE_Concat_input_pipe_39_inst_req_1); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_39_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Sample/rr
      -- 
    ca_158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_39_inst_ack_1, ack => concat_CP_34_elements(9)); -- 
    rr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(9), ack => type_cast_43_inst_req_0); -- 
    rr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(9), ack => RPIPE_Concat_input_pipe_51_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Sample/ra
      -- 
    ra_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_0, ack => concat_CP_34_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	76 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_43_Update/ca
      -- 
    ca_172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_1, ack => concat_CP_34_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_update_start_
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Update/cr
      -- 
    ra_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_51_inst_ack_0, ack => concat_CP_34_elements(12)); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(12), ack => RPIPE_Concat_input_pipe_51_inst_req_1); -- 
    -- CP-element group 13:  fork  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_51_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_51_inst_ack_1, ack => concat_CP_34_elements(13)); -- 
    rr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(13), ack => type_cast_55_inst_req_0); -- 
    rr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(13), ack => RPIPE_Concat_input_pipe_64_inst_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Sample/ra
      -- 
    ra_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_55_inst_ack_0, ack => concat_CP_34_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	76 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_55_Update/ca
      -- 
    ca_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_55_inst_ack_1, ack => concat_CP_34_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_update_start_
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Update/cr
      -- 
    ra_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_64_inst_ack_0, ack => concat_CP_34_elements(16)); -- 
    cr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(16), ack => RPIPE_Concat_input_pipe_64_inst_req_1); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	20 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_64_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Sample/rr
      -- 
    ca_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_64_inst_ack_1, ack => concat_CP_34_elements(17)); -- 
    rr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(17), ack => type_cast_68_inst_req_0); -- 
    rr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(17), ack => RPIPE_Concat_input_pipe_76_inst_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Sample/ra
      -- 
    ra_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_0, ack => concat_CP_34_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	76 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_68_Update/ca
      -- 
    ca_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_1, ack => concat_CP_34_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_update_start_
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Update/cr
      -- 
    ra_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_76_inst_ack_0, ack => concat_CP_34_elements(20)); -- 
    cr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(20), ack => RPIPE_Concat_input_pipe_76_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_76_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Sample/rr
      -- 
    ca_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_76_inst_ack_1, ack => concat_CP_34_elements(21)); -- 
    rr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(21), ack => type_cast_80_inst_req_0); -- 
    rr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(21), ack => RPIPE_Concat_input_pipe_89_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Sample/ra
      -- 
    ra_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_80_inst_ack_0, ack => concat_CP_34_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	76 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_80_Update/ca
      -- 
    ca_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_80_inst_ack_1, ack => concat_CP_34_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_update_start_
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Update/cr
      -- 
    ra_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_89_inst_ack_0, ack => concat_CP_34_elements(24)); -- 
    cr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(24), ack => RPIPE_Concat_input_pipe_89_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_89_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Sample/rr
      -- 
    ca_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_89_inst_ack_1, ack => concat_CP_34_elements(25)); -- 
    rr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(25), ack => type_cast_93_inst_req_0); -- 
    rr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(25), ack => RPIPE_Concat_input_pipe_101_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Sample/ra
      -- 
    ra_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_0, ack => concat_CP_34_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	76 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_93_Update/ca
      -- 
    ca_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_1, ack => concat_CP_34_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_update_start_
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Update/cr
      -- 
    ra_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_101_inst_ack_0, ack => concat_CP_34_elements(28)); -- 
    cr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(28), ack => RPIPE_Concat_input_pipe_101_inst_req_1); -- 
    -- CP-element group 29:  fork  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_101_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Sample/rr
      -- 
    ca_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_101_inst_ack_1, ack => concat_CP_34_elements(29)); -- 
    rr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(29), ack => type_cast_105_inst_req_0); -- 
    rr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(29), ack => RPIPE_Concat_input_pipe_114_inst_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Sample/ra
      -- 
    ra_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_0, ack => concat_CP_34_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	76 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_105_Update/ca
      -- 
    ca_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_1, ack => concat_CP_34_elements(31)); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	29 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_update_start_
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Update/cr
      -- 
    ra_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_114_inst_ack_0, ack => concat_CP_34_elements(32)); -- 
    cr_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(32), ack => RPIPE_Concat_input_pipe_114_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_114_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Sample/rr
      -- 
    ca_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_114_inst_ack_1, ack => concat_CP_34_elements(33)); -- 
    rr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(33), ack => RPIPE_Concat_input_pipe_126_inst_req_0); -- 
    rr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(33), ack => type_cast_118_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Sample/ra
      -- 
    ra_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_0, ack => concat_CP_34_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	0 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	76 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_118_Update/ca
      -- 
    ca_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_1, ack => concat_CP_34_elements(35)); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_update_start_
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Sample/ra
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Update/cr
      -- 
    ra_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_126_inst_ack_0, ack => concat_CP_34_elements(36)); -- 
    cr_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(36), ack => RPIPE_Concat_input_pipe_126_inst_req_1); -- 
    -- CP-element group 37:  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	40 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (9) 
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_126_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Sample/rr
      -- 
    ca_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_126_inst_ack_1, ack => concat_CP_34_elements(37)); -- 
    rr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(37), ack => type_cast_130_inst_req_0); -- 
    rr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(37), ack => RPIPE_Concat_input_pipe_139_inst_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Sample/ra
      -- 
    ra_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_0, ack => concat_CP_34_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	76 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_130_Update/ca
      -- 
    ca_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_1, ack => concat_CP_34_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Sample/ra
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Update/cr
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_update_start_
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Sample/$exit
      -- 
    ra_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_139_inst_ack_0, ack => concat_CP_34_elements(40)); -- 
    cr_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(40), ack => RPIPE_Concat_input_pipe_139_inst_req_1); -- 
    -- CP-element group 41:  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	44 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_139_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Sample/rr
      -- 
    ca_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_139_inst_ack_1, ack => concat_CP_34_elements(41)); -- 
    rr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(41), ack => RPIPE_Concat_input_pipe_151_inst_req_0); -- 
    rr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(41), ack => type_cast_143_inst_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Sample/ra
      -- 
    ra_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_0, ack => concat_CP_34_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	0 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	76 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_143_Update/ca
      -- 
    ca_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_1, ack => concat_CP_34_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	41 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_update_start_
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Update/cr
      -- 
    ra_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_151_inst_ack_0, ack => concat_CP_34_elements(44)); -- 
    cr_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(44), ack => RPIPE_Concat_input_pipe_151_inst_req_1); -- 
    -- CP-element group 45:  fork  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	48 
    -- CP-element group 45:  members (9) 
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_151_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Sample/rr
      -- 
    ca_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_151_inst_ack_1, ack => concat_CP_34_elements(45)); -- 
    rr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(45), ack => RPIPE_Concat_input_pipe_164_inst_req_0); -- 
    rr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(45), ack => type_cast_155_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Sample/ra
      -- 
    ra_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => concat_CP_34_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	76 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_155_Update/ca
      -- 
    ca_424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => concat_CP_34_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	45 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_update_start_
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Update/cr
      -- 
    ra_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_164_inst_ack_0, ack => concat_CP_34_elements(48)); -- 
    cr_437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(48), ack => RPIPE_Concat_input_pipe_164_inst_req_1); -- 
    -- CP-element group 49:  fork  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	52 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_164_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Sample/rr
      -- 
    ca_438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_164_inst_ack_1, ack => concat_CP_34_elements(49)); -- 
    rr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(49), ack => RPIPE_Concat_input_pipe_176_inst_req_0); -- 
    rr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(49), ack => type_cast_168_inst_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Sample/ra
      -- 
    ra_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_168_inst_ack_0, ack => concat_CP_34_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	0 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	76 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_168_Update/ca
      -- 
    ca_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_168_inst_ack_1, ack => concat_CP_34_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	49 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_update_start_
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Update/cr
      -- 
    ra_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_176_inst_ack_0, ack => concat_CP_34_elements(52)); -- 
    cr_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(52), ack => RPIPE_Concat_input_pipe_176_inst_req_1); -- 
    -- CP-element group 53:  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_176_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Sample/rr
      -- 
    ca_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_176_inst_ack_1, ack => concat_CP_34_elements(53)); -- 
    rr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(53), ack => type_cast_180_inst_req_0); -- 
    rr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(53), ack => RPIPE_Concat_input_pipe_189_inst_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Sample/ra
      -- 
    ra_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_180_inst_ack_0, ack => concat_CP_34_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	76 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_180_Update/ca
      -- 
    ca_480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_180_inst_ack_1, ack => concat_CP_34_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_update_start_
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Update/cr
      -- 
    ra_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_189_inst_ack_0, ack => concat_CP_34_elements(56)); -- 
    cr_493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(56), ack => RPIPE_Concat_input_pipe_189_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_189_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Sample/rr
      -- 
    ca_494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_189_inst_ack_1, ack => concat_CP_34_elements(57)); -- 
    rr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(57), ack => type_cast_193_inst_req_0); -- 
    rr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(57), ack => RPIPE_Concat_input_pipe_201_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Sample/ra
      -- 
    ra_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_0, ack => concat_CP_34_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	76 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_193_Update/ca
      -- 
    ca_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_1, ack => concat_CP_34_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	57 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_update_start_
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Sample/ra
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Update/cr
      -- 
    ra_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_201_inst_ack_0, ack => concat_CP_34_elements(60)); -- 
    cr_521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(60), ack => RPIPE_Concat_input_pipe_201_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: 	64 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_201_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Sample/rr
      -- 
    ca_522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_201_inst_ack_1, ack => concat_CP_34_elements(61)); -- 
    rr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(61), ack => type_cast_205_inst_req_0); -- 
    rr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(61), ack => RPIPE_Concat_input_pipe_214_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Sample/ra
      -- 
    ra_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_0, ack => concat_CP_34_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	0 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	76 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_205_Update/ca
      -- 
    ca_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_1, ack => concat_CP_34_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	61 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_update_start_
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Sample/ra
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Update/cr
      -- 
    ra_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_214_inst_ack_0, ack => concat_CP_34_elements(64)); -- 
    cr_549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(64), ack => RPIPE_Concat_input_pipe_214_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (9) 
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_214_Update/ca
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Sample/rr
      -- 
    ca_550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_214_inst_ack_1, ack => concat_CP_34_elements(65)); -- 
    rr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(65), ack => type_cast_218_inst_req_0); -- 
    rr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(65), ack => RPIPE_Concat_input_pipe_226_inst_req_0); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Sample/ra
      -- 
    ra_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_0, ack => concat_CP_34_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	76 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_218_Update/ca
      -- 
    ca_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_1, ack => concat_CP_34_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_update_start_
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Sample/ra
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Update/cr
      -- 
    ra_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_226_inst_ack_0, ack => concat_CP_34_elements(68)); -- 
    cr_577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(68), ack => RPIPE_Concat_input_pipe_226_inst_req_1); -- 
    -- CP-element group 69:  fork  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: 	72 
    -- CP-element group 69:  members (9) 
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_226_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Sample/rr
      -- 
    ca_578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_226_inst_ack_1, ack => concat_CP_34_elements(69)); -- 
    rr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(69), ack => type_cast_230_inst_req_0); -- 
    rr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(69), ack => RPIPE_Concat_input_pipe_239_inst_req_0); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Sample/ra
      -- 
    ra_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_230_inst_ack_0, ack => concat_CP_34_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	76 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_230_Update/ca
      -- 
    ca_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_230_inst_ack_1, ack => concat_CP_34_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	69 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_update_start_
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Update/cr
      -- 
    ra_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_239_inst_ack_0, ack => concat_CP_34_elements(72)); -- 
    cr_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(72), ack => RPIPE_Concat_input_pipe_239_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/RPIPE_Concat_input_pipe_239_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Sample/rr
      -- 
    ca_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_239_inst_ack_1, ack => concat_CP_34_elements(73)); -- 
    rr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(73), ack => type_cast_243_inst_req_0); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Sample/ra
      -- 
    ra_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_0, ack => concat_CP_34_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	0 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/type_cast_243_Update/ca
      -- 
    ca_620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_1, ack => concat_CP_34_elements(75)); -- 
    -- CP-element group 76:  branch  join  transition  place  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	63 
    -- CP-element group 76: 	55 
    -- CP-element group 76: 	51 
    -- CP-element group 76: 	59 
    -- CP-element group 76: 	39 
    -- CP-element group 76: 	43 
    -- CP-element group 76: 	35 
    -- CP-element group 76: 	47 
    -- CP-element group 76: 	67 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	75 
    -- CP-element group 76: 	7 
    -- CP-element group 76: 	11 
    -- CP-element group 76: 	15 
    -- CP-element group 76: 	19 
    -- CP-element group 76: 	23 
    -- CP-element group 76: 	27 
    -- CP-element group 76: 	31 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (10) 
      -- CP-element group 76: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297__exit__
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_298__entry__
      -- CP-element group 76: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_297/$exit
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_298_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_298_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_298_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_298_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_23/R_cmp467_299_place
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_298_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_298_else_link/$entry
      -- 
    branch_req_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(76), ack => if_stmt_298_branch_req_0); -- 
    concat_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 17) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1);
      constant place_markings: IntegerArray(0 to 17)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant place_delays: IntegerArray(0 to 17) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 18); -- 
    begin -- 
      preds <= concat_CP_34_elements(63) & concat_CP_34_elements(55) & concat_CP_34_elements(51) & concat_CP_34_elements(59) & concat_CP_34_elements(39) & concat_CP_34_elements(43) & concat_CP_34_elements(35) & concat_CP_34_elements(47) & concat_CP_34_elements(67) & concat_CP_34_elements(71) & concat_CP_34_elements(75) & concat_CP_34_elements(7) & concat_CP_34_elements(11) & concat_CP_34_elements(15) & concat_CP_34_elements(19) & concat_CP_34_elements(23) & concat_CP_34_elements(27) & concat_CP_34_elements(31);
      gj_concat_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 18, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: 	82 
    -- CP-element group 77:  members (18) 
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_319__exit__
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359__entry__
      -- CP-element group 77: 	 branch_block_stmt_23/if_stmt_298_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_23/if_stmt_298_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_23/entry_bbx_xnph469
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_update_start_
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_23/entry_bbx_xnph469_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/entry_bbx_xnph469_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_319_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_319_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_319_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_319_PhiAck/dummy
      -- 
    if_choice_transition_633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_298_branch_ack_1, ack => concat_CP_34_elements(77)); -- 
    rr_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(77), ack => type_cast_345_inst_req_0); -- 
    cr_677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(77), ack => type_cast_345_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	794 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_23/if_stmt_298_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_23/if_stmt_298_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_23/entry_forx_xcond163x_xpreheader
      -- CP-element group 78: 	 branch_block_stmt_23/entry_forx_xcond163x_xpreheader_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_23/entry_forx_xcond163x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_298_branch_ack_0, ack => concat_CP_34_elements(78)); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	794 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	194 
    -- CP-element group 79: 	195 
    -- CP-element group 79:  members (18) 
      -- CP-element group 79: 	 branch_block_stmt_23/merge_stmt_541__exit__
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581__entry__
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_update_start_
      -- CP-element group 79: 	 branch_block_stmt_23/if_stmt_313_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_23/if_stmt_313_if_link/if_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_23/forx_xcond163x_xpreheader_bbx_xnph465
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/$entry
      -- CP-element group 79: 	 branch_block_stmt_23/forx_xcond163x_xpreheader_bbx_xnph465_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_23/forx_xcond163x_xpreheader_bbx_xnph465_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_23/merge_stmt_541_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_23/merge_stmt_541_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_23/merge_stmt_541_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_23/merge_stmt_541_PhiAck/dummy
      -- 
    if_choice_transition_655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_313_branch_ack_1, ack => concat_CP_34_elements(79)); -- 
    cr_1106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(79), ack => type_cast_567_inst_req_1); -- 
    rr_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(79), ack => type_cast_567_inst_req_0); -- 
    -- CP-element group 80:  transition  place  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	794 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	795 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_23/if_stmt_313_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_23/if_stmt_313_else_link/else_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_23/forx_xcond163x_xpreheader_forx_xend223
      -- CP-element group 80: 	 branch_block_stmt_23/forx_xcond163x_xpreheader_forx_xend223_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_23/forx_xcond163x_xpreheader_forx_xend223_PhiReq/$exit
      -- 
    else_choice_transition_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_313_branch_ack_0, ack => concat_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Sample/ra
      -- 
    ra_673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => concat_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  place  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	77 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (13) 
      -- CP-element group 82: 	 branch_block_stmt_23/merge_stmt_361__exit__
      -- CP-element group 82: 	 branch_block_stmt_23/do_while_stmt_368__entry__
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359__exit__
      -- CP-element group 82: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/$exit
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_324_to_assign_stmt_359/type_cast_345_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/$entry
      -- CP-element group 82: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/$exit
      -- CP-element group 82: 	 branch_block_stmt_23/merge_stmt_361_PhiReqMerge
      -- CP-element group 82: 	 branch_block_stmt_23/merge_stmt_361_PhiAck/$entry
      -- CP-element group 82: 	 branch_block_stmt_23/merge_stmt_361_PhiAck/$exit
      -- 
    ca_678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => concat_CP_34_elements(82)); -- 
    -- CP-element group 83:  transition  place  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	89 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_23/do_while_stmt_368/$entry
      -- CP-element group 83: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368__entry__
      -- 
    concat_CP_34_elements(83) <= concat_CP_34_elements(82);
    -- CP-element group 84:  merge  place  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	191 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368__exit__
      -- 
    -- Element group concat_CP_34_elements(84) is bound as output of CP function.
    -- CP-element group 85:  merge  place  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	88 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_23/do_while_stmt_368/loop_back
      -- 
    -- Element group concat_CP_34_elements(85) is bound as output of CP function.
    -- CP-element group 86:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	91 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	189 
    -- CP-element group 86: 	190 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_23/do_while_stmt_368/loop_taken/$entry
      -- CP-element group 86: 	 branch_block_stmt_23/do_while_stmt_368/loop_exit/$entry
      -- CP-element group 86: 	 branch_block_stmt_23/do_while_stmt_368/condition_done
      -- 
    concat_CP_34_elements(86) <= concat_CP_34_elements(91);
    -- CP-element group 87:  branch  place  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	188 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_23/do_while_stmt_368/loop_body_done
      -- 
    concat_CP_34_elements(87) <= concat_CP_34_elements(188);
    -- CP-element group 88:  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	85 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	97 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/back_edge_to_loop_body
      -- 
    concat_CP_34_elements(88) <= concat_CP_34_elements(85);
    -- CP-element group 89:  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	83 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	99 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/first_time_through_loop_body
      -- 
    concat_CP_34_elements(89) <= concat_CP_34_elements(83);
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	93 
    -- CP-element group 90: 	94 
    -- CP-element group 90: 	113 
    -- CP-element group 90: 	114 
    -- CP-element group 90: 	119 
    -- CP-element group 90: 	187 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/$entry
      -- CP-element group 90: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/loop_body_start
      -- 
    -- Element group concat_CP_34_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	96 
    -- CP-element group 91: 	187 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	86 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/condition_evaluated
      -- 
    condition_evaluated_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(91), ack => do_while_stmt_368_branch_req_0); -- 
    concat_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(96) & concat_CP_34_elements(187);
      gj_concat_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	96 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/aggregated_phi_sample_req
      -- CP-element group 92: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_sample_start__ps
      -- 
    concat_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(93) & concat_CP_34_elements(96);
      gj_concat_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	92 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_sample_start_
      -- 
    concat_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 26) := "concat_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(90) & concat_CP_34_elements(95);
      gj_concat_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	90 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: 	115 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/aggregated_phi_update_req
      -- CP-element group 94: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_update_start_
      -- CP-element group 94: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_update_start__ps
      -- 
    concat_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 26) := "concat_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(90) & concat_CP_34_elements(96) & concat_CP_34_elements(115);
      gj_concat_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	188 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/aggregated_phi_sample_ack
      -- CP-element group 95: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(95) is bound as output of CP function.
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	91 
    -- CP-element group 96: 	115 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (16) 
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_resized_1
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_scaled_1
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_computed_1
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_resize_1/$entry
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_resize_1/$exit
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_resize_1/index_resize_req
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_resize_1/index_resize_ack
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_scale_1/$entry
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_scale_1/$exit
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_scale_1/scale_rename_req
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_index_scale_1/scale_rename_ack
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/aggregated_phi_update_ack
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Sample/req
      -- 
    req_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(96), ack => array_obj_ref_380_index_offset_req_0); -- 
    -- Element group concat_CP_34_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	88 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_loopback_trigger
      -- 
    concat_CP_34_elements(97) <= concat_CP_34_elements(88);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_loopback_sample_req
      -- CP-element group 98: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_loopback_sample_req_ps
      -- 
    phi_stmt_370_loopback_sample_req_708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_370_loopback_sample_req_708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(98), ack => phi_stmt_370_req_0); -- 
    -- Element group concat_CP_34_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	89 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_entry_trigger
      -- 
    concat_CP_34_elements(99) <= concat_CP_34_elements(89);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_entry_sample_req
      -- CP-element group 100: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_entry_sample_req_ps
      -- 
    phi_stmt_370_entry_sample_req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_370_entry_sample_req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(100), ack => phi_stmt_370_req_1); -- 
    -- Element group concat_CP_34_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_phi_mux_ack
      -- CP-element group 101: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/phi_stmt_370_phi_mux_ack_ps
      -- 
    phi_stmt_370_phi_mux_ack_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_370_ack_0, ack => concat_CP_34_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Sample/rr
      -- 
    rr_727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(104), ack => type_cast_373_inst_req_0); -- 
    concat_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(102) & concat_CP_34_elements(106);
      gj_concat_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_update_start_
      -- CP-element group 105: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Update/cr
      -- 
    cr_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(105), ack => type_cast_373_inst_req_1); -- 
    concat_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(103) & concat_CP_34_elements(107);
      gj_concat_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Sample/ra
      -- 
    ra_728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_373_inst_ack_0, ack => concat_CP_34_elements(106)); -- 
    -- CP-element group 107:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_373_Update/ca
      -- 
    ca_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_373_inst_ack_1, ack => concat_CP_34_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_sample_start__ps
      -- CP-element group 108: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_update_start__ps
      -- CP-element group 109: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_update_start_
      -- 
    -- Element group concat_CP_34_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_update_completed__ps
      -- 
    concat_CP_34_elements(110) <= concat_CP_34_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/R_indvar488_at_entry_374_update_completed_
      -- 
    -- Element group concat_CP_34_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => concat_CP_34_elements(109), ack => concat_CP_34_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	116 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	117 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	117 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_request/$entry
      -- CP-element group 112: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_request/req
      -- 
    req_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(112), ack => addr_of_381_final_reg_req_0); -- 
    concat_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(116) & concat_CP_34_elements(117);
      gj_concat_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	90 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	118 
    -- CP-element group 113: 	185 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_update_start_
      -- CP-element group 113: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_complete/$entry
      -- CP-element group 113: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_complete/req
      -- 
    req_787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(113), ack => addr_of_381_final_reg_req_1); -- 
    concat_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(90) & concat_CP_34_elements(118) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	90 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: 	117 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_update_start
      -- CP-element group 114: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Update/req
      -- 
    req_772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(114), ack => array_obj_ref_380_index_offset_req_1); -- 
    concat_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(90) & concat_CP_34_elements(116) & concat_CP_34_elements(117);
      gj_concat_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	96 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	188 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	94 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_sample_complete
      -- CP-element group 115: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Sample/ack
      -- 
    ack_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_380_index_offset_ack_0, ack => concat_CP_34_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	112 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (8) 
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_offset_calculated
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_final_index_sum_regn_Update/ack
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_base_plus_offset/$entry
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_base_plus_offset/$exit
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_base_plus_offset/sum_rename_req
      -- CP-element group 116: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/array_obj_ref_380_base_plus_offset/sum_rename_ack
      -- 
    ack_773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_380_index_offset_ack_1, ack => concat_CP_34_elements(116)); -- 
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	112 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	112 
    -- CP-element group 117: 	114 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_request/$exit
      -- CP-element group 117: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_request/ack
      -- 
    ack_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_381_final_reg_ack_0, ack => concat_CP_34_elements(117)); -- 
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	113 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	183 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	113 
    -- CP-element group 118:  members (19) 
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_root_address_calculated
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_word_address_calculated
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_address_calculated
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_word_addrgen/root_register_ack
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_word_addrgen/root_register_req
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_word_addrgen/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_word_addrgen/$entry
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_plus_offset/sum_rename_ack
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_plus_offset/sum_rename_req
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_plus_offset/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_plus_offset/$entry
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_addr_resize/base_resize_ack
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_addr_resize/base_resize_req
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_addr_resize/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_addr_resize/$entry
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_base_address_resized
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/addr_of_381_complete/ack
      -- 
    ack_788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_381_final_reg_ack_1, ack => concat_CP_34_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	90 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	122 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Sample/rr
      -- 
    rr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(119), ack => RPIPE_Concat_input_pipe_384_inst_req_0); -- 
    concat_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(90) & concat_CP_34_elements(122);
      gj_concat_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	125 
    -- CP-element group 120: 	178 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_update_start_
      -- CP-element group 120: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Update/cr
      -- 
    cr_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(120), ack => RPIPE_Concat_input_pipe_384_inst_req_1); -- 
    concat_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(121) & concat_CP_34_elements(125) & concat_CP_34_elements(178);
      gj_concat_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	120 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Sample/ra
      -- 
    ra_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_384_inst_ack_0, ack => concat_CP_34_elements(121)); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122: 	127 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	119 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_384_Update/ca
      -- 
    ca_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_384_inst_ack_1, ack => concat_CP_34_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Sample/rr
      -- 
    rr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(123), ack => type_cast_388_inst_req_0); -- 
    concat_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(122) & concat_CP_34_elements(125);
      gj_concat_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: 	185 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_update_start_
      -- CP-element group 124: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Update/cr
      -- 
    cr_815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(124), ack => type_cast_388_inst_req_1); -- 
    concat_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(126) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	120 
    -- CP-element group 125: 	123 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Sample/ra
      -- 
    ra_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_388_inst_ack_0, ack => concat_CP_34_elements(125)); -- 
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	183 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_388_Update/ca
      -- 
    ca_816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_388_inst_ack_1, ack => concat_CP_34_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	122 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	130 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Sample/rr
      -- 
    rr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(127), ack => RPIPE_Concat_input_pipe_397_inst_req_0); -- 
    concat_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(122) & concat_CP_34_elements(130);
      gj_concat_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	129 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_update_start_
      -- CP-element group 128: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Update/cr
      -- 
    cr_829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(128), ack => RPIPE_Concat_input_pipe_397_inst_req_1); -- 
    concat_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(129) & concat_CP_34_elements(133);
      gj_concat_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	128 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Sample/ra
      -- 
    ra_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_397_inst_ack_0, ack => concat_CP_34_elements(129)); -- 
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	135 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	127 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_397_Update/ca
      -- 
    ca_830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_397_inst_ack_1, ack => concat_CP_34_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Sample/rr
      -- 
    rr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(131), ack => type_cast_401_inst_req_0); -- 
    concat_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(130) & concat_CP_34_elements(133);
      gj_concat_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	185 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_update_start_
      -- CP-element group 132: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Update/cr
      -- 
    cr_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(132), ack => type_cast_401_inst_req_1); -- 
    concat_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(134) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Sample/ra
      -- 
    ra_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_401_inst_ack_0, ack => concat_CP_34_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	183 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_401_Update/ca
      -- 
    ca_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_401_inst_ack_1, ack => concat_CP_34_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	130 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	138 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Sample/rr
      -- 
    rr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(135), ack => RPIPE_Concat_input_pipe_415_inst_req_0); -- 
    concat_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(130) & concat_CP_34_elements(138);
      gj_concat_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	137 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	141 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_update_start_
      -- CP-element group 136: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Update/cr
      -- 
    cr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(136), ack => RPIPE_Concat_input_pipe_415_inst_req_1); -- 
    concat_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(137) & concat_CP_34_elements(141);
      gj_concat_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	136 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Sample/ra
      -- 
    ra_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_415_inst_ack_0, ack => concat_CP_34_elements(137)); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	143 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	135 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_415_Update/ca
      -- 
    ca_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_415_inst_ack_1, ack => concat_CP_34_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Sample/rr
      -- 
    rr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(139), ack => type_cast_419_inst_req_0); -- 
    concat_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(138) & concat_CP_34_elements(141);
      gj_concat_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: 	185 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_update_start_
      -- CP-element group 140: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Update/cr
      -- 
    cr_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(140), ack => type_cast_419_inst_req_1); -- 
    concat_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(142) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	136 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Sample/ra
      -- 
    ra_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_419_inst_ack_0, ack => concat_CP_34_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	183 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_419_Update/ca
      -- 
    ca_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_419_inst_ack_1, ack => concat_CP_34_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	138 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	146 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Sample/rr
      -- 
    rr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(143), ack => RPIPE_Concat_input_pipe_433_inst_req_0); -- 
    concat_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(138) & concat_CP_34_elements(146);
      gj_concat_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	145 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	149 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_update_start_
      -- CP-element group 144: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Update/cr
      -- 
    cr_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(144), ack => RPIPE_Concat_input_pipe_433_inst_req_1); -- 
    concat_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(145) & concat_CP_34_elements(149);
      gj_concat_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	144 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Sample/ra
      -- 
    ra_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_433_inst_ack_0, ack => concat_CP_34_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	151 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	143 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_433_Update/ca
      -- 
    ca_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_433_inst_ack_1, ack => concat_CP_34_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Sample/rr
      -- 
    rr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(147), ack => type_cast_437_inst_req_0); -- 
    concat_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(146) & concat_CP_34_elements(149);
      gj_concat_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: 	185 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_update_start_
      -- CP-element group 148: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Update/cr
      -- 
    cr_899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(148), ack => type_cast_437_inst_req_1); -- 
    concat_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(150) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	144 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Sample/ra
      -- 
    ra_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_437_inst_ack_0, ack => concat_CP_34_elements(149)); -- 
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	183 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_437_Update/ca
      -- 
    ca_900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_437_inst_ack_1, ack => concat_CP_34_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	146 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	154 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Sample/rr
      -- 
    rr_908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(151), ack => RPIPE_Concat_input_pipe_451_inst_req_0); -- 
    concat_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(146) & concat_CP_34_elements(154);
      gj_concat_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	153 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	157 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_update_start_
      -- CP-element group 152: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Update/cr
      -- 
    cr_913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(152), ack => RPIPE_Concat_input_pipe_451_inst_req_1); -- 
    concat_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(153) & concat_CP_34_elements(157);
      gj_concat_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	152 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Sample/ra
      -- 
    ra_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_451_inst_ack_0, ack => concat_CP_34_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	159 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	151 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_451_Update/ca
      -- 
    ca_914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_451_inst_ack_1, ack => concat_CP_34_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Sample/rr
      -- 
    rr_922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(155), ack => type_cast_455_inst_req_0); -- 
    concat_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(154) & concat_CP_34_elements(157);
      gj_concat_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: 	185 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_update_start_
      -- CP-element group 156: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Update/cr
      -- 
    cr_927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(156), ack => type_cast_455_inst_req_1); -- 
    concat_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(158) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	152 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Sample/ra
      -- 
    ra_923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_455_inst_ack_0, ack => concat_CP_34_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	183 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_455_Update/ca
      -- 
    ca_928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_455_inst_ack_1, ack => concat_CP_34_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	154 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	162 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Sample/rr
      -- 
    rr_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(159), ack => RPIPE_Concat_input_pipe_469_inst_req_0); -- 
    concat_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(154) & concat_CP_34_elements(162);
      gj_concat_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	161 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	165 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_update_start_
      -- CP-element group 160: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Update/cr
      -- 
    cr_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(160), ack => RPIPE_Concat_input_pipe_469_inst_req_1); -- 
    concat_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(161) & concat_CP_34_elements(165);
      gj_concat_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	160 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Sample/ra
      -- 
    ra_937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_469_inst_ack_0, ack => concat_CP_34_elements(161)); -- 
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	167 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	159 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_469_Update/ca
      -- 
    ca_942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_469_inst_ack_1, ack => concat_CP_34_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_sample_start_
      -- 
    rr_950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(163), ack => type_cast_473_inst_req_0); -- 
    concat_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(162) & concat_CP_34_elements(165);
      gj_concat_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: 	185 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Update/cr
      -- CP-element group 164: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_update_start_
      -- 
    cr_955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(164), ack => type_cast_473_inst_req_1); -- 
    concat_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(166) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	160 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Sample/ra
      -- CP-element group 165: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_sample_completed_
      -- 
    ra_951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_0, ack => concat_CP_34_elements(165)); -- 
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	183 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_473_update_completed_
      -- 
    ca_956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_1, ack => concat_CP_34_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	162 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	170 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Sample/$entry
      -- 
    rr_964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(167), ack => RPIPE_Concat_input_pipe_487_inst_req_0); -- 
    concat_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(162) & concat_CP_34_elements(170);
      gj_concat_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	173 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_update_start_
      -- 
    cr_969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(168), ack => RPIPE_Concat_input_pipe_487_inst_req_1); -- 
    concat_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(169) & concat_CP_34_elements(173);
      gj_concat_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	168 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Sample/ra
      -- CP-element group 169: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_sample_completed_
      -- 
    ra_965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_487_inst_ack_0, ack => concat_CP_34_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170: 	175 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	167 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_Update/ca
      -- CP-element group 170: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_487_update_completed_
      -- 
    ca_970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_487_inst_ack_1, ack => concat_CP_34_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Sample/rr
      -- CP-element group 171: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Sample/$entry
      -- 
    rr_978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(171), ack => type_cast_491_inst_req_0); -- 
    concat_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(170) & concat_CP_34_elements(173);
      gj_concat_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: 	185 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_update_start_
      -- CP-element group 172: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Update/$entry
      -- 
    cr_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(172), ack => type_cast_491_inst_req_1); -- 
    concat_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(174) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	168 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Sample/$exit
      -- 
    ra_979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_0, ack => concat_CP_34_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	183 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_491_Update/$exit
      -- 
    ca_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_1, ack => concat_CP_34_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	170 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	178 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_sample_start_
      -- 
    rr_992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(175), ack => RPIPE_Concat_input_pipe_505_inst_req_0); -- 
    concat_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(170) & concat_CP_34_elements(178);
      gj_concat_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	181 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Update/cr
      -- CP-element group 176: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_update_start_
      -- 
    cr_997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(176), ack => RPIPE_Concat_input_pipe_505_inst_req_1); -- 
    concat_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(177) & concat_CP_34_elements(181);
      gj_concat_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	176 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Sample/$exit
      -- 
    ra_993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_505_inst_ack_0, ack => concat_CP_34_elements(177)); -- 
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	120 
    -- CP-element group 178: 	175 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/RPIPE_Concat_input_pipe_505_update_completed_
      -- 
    ca_998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_505_inst_ack_1, ack => concat_CP_34_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Sample/rr
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_sample_start_
      -- 
    rr_1006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(179), ack => type_cast_509_inst_req_0); -- 
    concat_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(178) & concat_CP_34_elements(181);
      gj_concat_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: 	185 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Update/cr
      -- CP-element group 180: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_update_start_
      -- 
    cr_1011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(180), ack => type_cast_509_inst_req_1); -- 
    concat_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(182) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	176 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_sample_completed_
      -- 
    ra_1007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_509_inst_ack_0, ack => concat_CP_34_elements(181)); -- 
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/type_cast_509_Update/$exit
      -- 
    ca_1012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_509_inst_ack_1, ack => concat_CP_34_elements(182)); -- 
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	118 
    -- CP-element group 183: 	126 
    -- CP-element group 183: 	134 
    -- CP-element group 183: 	142 
    -- CP-element group 183: 	150 
    -- CP-element group 183: 	158 
    -- CP-element group 183: 	166 
    -- CP-element group 183: 	174 
    -- CP-element group 183: 	182 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (9) 
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/word_access_start/word_0/rr
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/word_access_start/word_0/$entry
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/word_access_start/$entry
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/ptr_deref_517_Split/split_ack
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/ptr_deref_517_Split/split_req
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/ptr_deref_517_Split/$exit
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/ptr_deref_517_Split/$entry
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/$entry
      -- 
    rr_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(183), ack => ptr_deref_517_store_0_req_0); -- 
    concat_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= concat_CP_34_elements(118) & concat_CP_34_elements(126) & concat_CP_34_elements(134) & concat_CP_34_elements(142) & concat_CP_34_elements(150) & concat_CP_34_elements(158) & concat_CP_34_elements(166) & concat_CP_34_elements(174) & concat_CP_34_elements(182) & concat_CP_34_elements(185);
      gj_concat_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (5) 
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_update_start_
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/word_access_complete/word_0/cr
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/word_access_complete/word_0/$entry
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/word_access_complete/$entry
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/$entry
      -- 
    cr_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(184), ack => ptr_deref_517_store_0_req_1); -- 
    concat_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(186);
      gj_concat_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	113 
    -- CP-element group 185: 	124 
    -- CP-element group 185: 	132 
    -- CP-element group 185: 	140 
    -- CP-element group 185: 	148 
    -- CP-element group 185: 	156 
    -- CP-element group 185: 	164 
    -- CP-element group 185: 	172 
    -- CP-element group 185: 	180 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (5) 
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/word_access_start/word_0/ra
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/word_access_start/word_0/$exit
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/word_access_start/$exit
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Sample/$exit
      -- 
    ra_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_517_store_0_ack_0, ack => concat_CP_34_elements(185)); -- 
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (5) 
      -- CP-element group 186: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/word_access_complete/word_0/ca
      -- CP-element group 186: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/word_access_complete/word_0/$exit
      -- CP-element group 186: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/word_access_complete/$exit
      -- CP-element group 186: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/ptr_deref_517_Update/$exit
      -- 
    ca_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_517_store_0_ack_1, ack => concat_CP_34_elements(186)); -- 
    -- CP-element group 187:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	90 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	91 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group concat_CP_34_elements(187) is a control-delay.
    cp_element_187_delay: control_delay_element  generic map(name => " 187_delay", delay_value => 1)  port map(req => concat_CP_34_elements(90), ack => concat_CP_34_elements(187), clk => clk, reset =>reset);
    -- CP-element group 188:  join  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	95 
    -- CP-element group 188: 	115 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	87 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_23/do_while_stmt_368/do_while_stmt_368_loop_body/$exit
      -- 
    concat_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(95) & concat_CP_34_elements(115) & concat_CP_34_elements(186);
      gj_concat_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	86 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_23/do_while_stmt_368/loop_exit/ack
      -- CP-element group 189: 	 branch_block_stmt_23/do_while_stmt_368/loop_exit/$exit
      -- 
    ack_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_368_branch_ack_0, ack => concat_CP_34_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	86 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_23/do_while_stmt_368/loop_taken/ack
      -- CP-element group 190: 	 branch_block_stmt_23/do_while_stmt_368/loop_taken/$exit
      -- 
    ack_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_368_branch_ack_1, ack => concat_CP_34_elements(190)); -- 
    -- CP-element group 191:  transition  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	84 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	1 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 branch_block_stmt_23/do_while_stmt_368/$exit
      -- 
    concat_CP_34_elements(191) <= concat_CP_34_elements(84);
    -- CP-element group 192:  merge  transition  place  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	1 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	794 
    -- CP-element group 192:  members (13) 
      -- CP-element group 192: 	 branch_block_stmt_23/if_stmt_537_if_link/if_choice_transition
      -- CP-element group 192: 	 branch_block_stmt_23/merge_stmt_304__exit__
      -- CP-element group 192: 	 branch_block_stmt_23/forx_xcond163x_xpreheaderx_xloopexit_forx_xcond163x_xpreheader
      -- CP-element group 192: 	 branch_block_stmt_23/if_stmt_537_if_link/$exit
      -- CP-element group 192: 	 branch_block_stmt_23/forx_xbody_forx_xcond163x_xpreheaderx_xloopexit
      -- CP-element group 192: 	 branch_block_stmt_23/forx_xbody_forx_xcond163x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 192: 	 branch_block_stmt_23/forx_xbody_forx_xcond163x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 192: 	 branch_block_stmt_23/merge_stmt_304_PhiReqMerge
      -- CP-element group 192: 	 branch_block_stmt_23/merge_stmt_304_PhiAck/$entry
      -- CP-element group 192: 	 branch_block_stmt_23/merge_stmt_304_PhiAck/$exit
      -- CP-element group 192: 	 branch_block_stmt_23/merge_stmt_304_PhiAck/dummy
      -- CP-element group 192: 	 branch_block_stmt_23/forx_xcond163x_xpreheaderx_xloopexit_forx_xcond163x_xpreheader_PhiReq/$entry
      -- CP-element group 192: 	 branch_block_stmt_23/forx_xcond163x_xpreheaderx_xloopexit_forx_xcond163x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_537_branch_ack_1, ack => concat_CP_34_elements(192)); -- 
    -- CP-element group 193:  merge  transition  place  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	1 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (5) 
      -- CP-element group 193: 	 branch_block_stmt_23/if_stmt_537_else_link/$exit
      -- CP-element group 193: 	 branch_block_stmt_23/if_stmt_537__exit__
      -- CP-element group 193: 	 branch_block_stmt_23/merge_stmt_541__entry__
      -- CP-element group 193: 	 branch_block_stmt_23/if_stmt_537_else_link/else_choice_transition
      -- CP-element group 193: 	 branch_block_stmt_23/merge_stmt_541_dead_link/$entry
      -- 
    else_choice_transition_1089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_537_branch_ack_0, ack => concat_CP_34_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	79 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_sample_completed_
      -- 
    ra_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_567_inst_ack_0, ack => concat_CP_34_elements(194)); -- 
    -- CP-element group 195:  transition  place  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	79 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (13) 
      -- CP-element group 195: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581__exit__
      -- CP-element group 195: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody169
      -- CP-element group 195: 	 branch_block_stmt_23/merge_stmt_583__exit__
      -- CP-element group 195: 	 branch_block_stmt_23/do_while_stmt_590__entry__
      -- CP-element group 195: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/type_cast_567_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_23/assign_stmt_546_to_assign_stmt_581/$exit
      -- CP-element group 195: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody169_PhiReq/$entry
      -- CP-element group 195: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody169_PhiReq/$exit
      -- CP-element group 195: 	 branch_block_stmt_23/merge_stmt_583_PhiReqMerge
      -- CP-element group 195: 	 branch_block_stmt_23/merge_stmt_583_PhiAck/$entry
      -- CP-element group 195: 	 branch_block_stmt_23/merge_stmt_583_PhiAck/$exit
      -- 
    ca_1107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_567_inst_ack_1, ack => concat_CP_34_elements(195)); -- 
    -- CP-element group 196:  transition  place  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	202 
    -- CP-element group 196:  members (2) 
      -- CP-element group 196: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590__entry__
      -- CP-element group 196: 	 branch_block_stmt_23/do_while_stmt_590/$entry
      -- 
    concat_CP_34_elements(196) <= concat_CP_34_elements(195);
    -- CP-element group 197:  merge  place  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	304 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590__exit__
      -- 
    -- Element group concat_CP_34_elements(197) is bound as output of CP function.
    -- CP-element group 198:  merge  place  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_23/do_while_stmt_590/loop_back
      -- 
    -- Element group concat_CP_34_elements(198) is bound as output of CP function.
    -- CP-element group 199:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	204 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	302 
    -- CP-element group 199: 	303 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_23/do_while_stmt_590/condition_done
      -- CP-element group 199: 	 branch_block_stmt_23/do_while_stmt_590/loop_exit/$entry
      -- CP-element group 199: 	 branch_block_stmt_23/do_while_stmt_590/loop_taken/$entry
      -- 
    concat_CP_34_elements(199) <= concat_CP_34_elements(204);
    -- CP-element group 200:  branch  place  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	301 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_23/do_while_stmt_590/loop_body_done
      -- 
    concat_CP_34_elements(200) <= concat_CP_34_elements(301);
    -- CP-element group 201:  transition  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	210 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/back_edge_to_loop_body
      -- 
    concat_CP_34_elements(201) <= concat_CP_34_elements(198);
    -- CP-element group 202:  transition  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	196 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	212 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/first_time_through_loop_body
      -- 
    concat_CP_34_elements(202) <= concat_CP_34_elements(196);
    -- CP-element group 203:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	206 
    -- CP-element group 203: 	207 
    -- CP-element group 203: 	226 
    -- CP-element group 203: 	227 
    -- CP-element group 203: 	232 
    -- CP-element group 203: 	300 
    -- CP-element group 203:  members (2) 
      -- CP-element group 203: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/$entry
      -- CP-element group 203: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/loop_body_start
      -- 
    -- Element group concat_CP_34_elements(203) is bound as output of CP function.
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	209 
    -- CP-element group 204: 	300 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	199 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/condition_evaluated
      -- 
    condition_evaluated_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(204), ack => do_while_stmt_590_branch_req_0); -- 
    concat_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(209) & concat_CP_34_elements(300);
      gj_concat_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	206 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	209 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_sample_start__ps
      -- CP-element group 205: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/aggregated_phi_sample_req
      -- 
    concat_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(206) & concat_CP_34_elements(209);
      gj_concat_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  join  transition  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	203 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	205 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_sample_start_
      -- 
    concat_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(203) & concat_CP_34_elements(208);
      gj_concat_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	203 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: 	228 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_update_start__ps
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_update_start_
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/aggregated_phi_update_req
      -- 
    concat_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(203) & concat_CP_34_elements(209) & concat_CP_34_elements(228);
      gj_concat_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	301 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_sample_completed__ps
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/aggregated_phi_sample_ack
      -- 
    -- Element group concat_CP_34_elements(208) is bound as output of CP function.
    -- CP-element group 209:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	204 
    -- CP-element group 209: 	228 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	205 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (16) 
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_resize_1/index_resize_req
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_resize_1/$exit
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_resize_1/$entry
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_computed_1
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_scaled_1
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_resized_1
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_update_completed__ps
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Sample/req
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Sample/$entry
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/aggregated_phi_update_ack
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_scale_1/scale_rename_ack
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_scale_1/scale_rename_req
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_scale_1/$exit
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_scale_1/$entry
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_index_resize_1/index_resize_ack
      -- 
    req_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(209), ack => array_obj_ref_602_index_offset_req_0); -- 
    -- Element group concat_CP_34_elements(209) is bound as output of CP function.
    -- CP-element group 210:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	201 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_loopback_trigger
      -- 
    concat_CP_34_elements(210) <= concat_CP_34_elements(201);
    -- CP-element group 211:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (2) 
      -- CP-element group 211: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_loopback_sample_req_ps
      -- CP-element group 211: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_loopback_sample_req
      -- 
    phi_stmt_592_loopback_sample_req_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_592_loopback_sample_req_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(211), ack => phi_stmt_592_req_0); -- 
    -- Element group concat_CP_34_elements(211) is bound as output of CP function.
    -- CP-element group 212:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	202 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_entry_trigger
      -- 
    concat_CP_34_elements(212) <= concat_CP_34_elements(202);
    -- CP-element group 213:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (2) 
      -- CP-element group 213: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_entry_sample_req_ps
      -- CP-element group 213: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_entry_sample_req
      -- 
    phi_stmt_592_entry_sample_req_1140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_592_entry_sample_req_1140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(213), ack => phi_stmt_592_req_1); -- 
    -- Element group concat_CP_34_elements(213) is bound as output of CP function.
    -- CP-element group 214:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (2) 
      -- CP-element group 214: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_phi_mux_ack_ps
      -- CP-element group 214: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/phi_stmt_592_phi_mux_ack
      -- 
    phi_stmt_592_phi_mux_ack_1143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_592_ack_0, ack => concat_CP_34_elements(214)); -- 
    -- CP-element group 215:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(215) is bound as output of CP function.
    -- CP-element group 216:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (1) 
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(216) is bound as output of CP function.
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Sample/rr
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_sample_start_
      -- 
    rr_1156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(217), ack => type_cast_595_inst_req_0); -- 
    concat_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(215) & concat_CP_34_elements(219);
      gj_concat_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_update_start_
      -- 
    cr_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(218), ack => type_cast_595_inst_req_1); -- 
    concat_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(216) & concat_CP_34_elements(220);
      gj_concat_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (4) 
      -- CP-element group 219: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Sample/ra
      -- CP-element group 219: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_sample_completed__ps
      -- 
    ra_1157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_0, ack => concat_CP_34_elements(219)); -- 
    -- CP-element group 220:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	218 
    -- CP-element group 220:  members (4) 
      -- CP-element group 220: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Update/ca
      -- CP-element group 220: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_595_update_completed__ps
      -- 
    ca_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_1, ack => concat_CP_34_elements(220)); -- 
    -- CP-element group 221:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (4) 
      -- CP-element group 221: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_sample_completed__ps
      -- CP-element group 221: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(221) is bound as output of CP function.
    -- CP-element group 222:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (2) 
      -- CP-element group 222: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_update_start_
      -- CP-element group 222: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(222) is bound as output of CP function.
    -- CP-element group 223:  join  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_update_completed__ps
      -- 
    concat_CP_34_elements(223) <= concat_CP_34_elements(224);
    -- CP-element group 224:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	223 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/R_indvar476_at_entry_596_update_completed_
      -- 
    -- Element group concat_CP_34_elements(224) is a control-delay.
    cp_element_224_delay: control_delay_element  generic map(name => " 224_delay", delay_value => 1)  port map(req => concat_CP_34_elements(222), ack => concat_CP_34_elements(224), clk => clk, reset =>reset);
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	229 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	230 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	230 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_request/$entry
      -- CP-element group 225: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_request/req
      -- 
    req_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(225), ack => addr_of_603_final_reg_req_0); -- 
    concat_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(229) & concat_CP_34_elements(230);
      gj_concat_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	203 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	231 
    -- CP-element group 226: 	298 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	231 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_update_start_
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_complete/req
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_complete/$entry
      -- 
    req_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(226), ack => addr_of_603_final_reg_req_1); -- 
    concat_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(203) & concat_CP_34_elements(231) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	203 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	229 
    -- CP-element group 227: 	230 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Update/req
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_update_start
      -- 
    req_1201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(227), ack => array_obj_ref_602_index_offset_req_1); -- 
    concat_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(203) & concat_CP_34_elements(229) & concat_CP_34_elements(230);
      gj_concat_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	209 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	301 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	207 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Sample/ack
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_sample_complete
      -- 
    ack_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_602_index_offset_ack_0, ack => concat_CP_34_elements(228)); -- 
    -- CP-element group 229:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	225 
    -- CP-element group 229: marked-successors 
    -- CP-element group 229: 	227 
    -- CP-element group 229:  members (8) 
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_base_plus_offset/$entry
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_offset_calculated
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_root_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_base_plus_offset/sum_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_base_plus_offset/sum_rename_req
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Update/ack
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_base_plus_offset/$exit
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/array_obj_ref_602_final_index_sum_regn_Update/$exit
      -- 
    ack_1202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_602_index_offset_ack_1, ack => concat_CP_34_elements(229)); -- 
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	225 
    -- CP-element group 230: successors 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	225 
    -- CP-element group 230: 	227 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_request/ack
      -- CP-element group 230: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_request/$exit
      -- 
    ack_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_603_final_reg_ack_0, ack => concat_CP_34_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	226 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	296 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	226 
    -- CP-element group 231:  members (19) 
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_complete/ack
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/addr_of_603_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_address_calculated
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_word_address_calculated
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_root_address_calculated
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_address_resized
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_addr_resize/$entry
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_addr_resize/$exit
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_addr_resize/base_resize_req
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_addr_resize/base_resize_ack
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_plus_offset/$entry
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_plus_offset/$exit
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_plus_offset/sum_rename_req
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_base_plus_offset/sum_rename_ack
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_word_addrgen/$entry
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_word_addrgen/$exit
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_word_addrgen/root_register_req
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_word_addrgen/root_register_ack
      -- 
    ack_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_603_final_reg_ack_1, ack => concat_CP_34_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	203 
    -- CP-element group 232: marked-predecessors 
    -- CP-element group 232: 	235 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Sample/rr
      -- CP-element group 232: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_sample_start_
      -- 
    rr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(232), ack => RPIPE_Concat_input_pipe_606_inst_req_0); -- 
    concat_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(203) & concat_CP_34_elements(235);
      gj_concat_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	234 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	238 
    -- CP-element group 233: 	291 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_update_start_
      -- 
    cr_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(233), ack => RPIPE_Concat_input_pipe_606_inst_req_1); -- 
    concat_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(234) & concat_CP_34_elements(238) & concat_CP_34_elements(291);
      gj_concat_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  transition  input  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	233 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Sample/ra
      -- CP-element group 234: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_sample_completed_
      -- 
    ra_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_606_inst_ack_0, ack => concat_CP_34_elements(234)); -- 
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235: 	240 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	232 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Update/ca
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_606_update_completed_
      -- 
    ca_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_606_inst_ack_1, ack => concat_CP_34_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: marked-predecessors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Sample/rr
      -- CP-element group 236: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_sample_start_
      -- 
    rr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(236), ack => type_cast_610_inst_req_0); -- 
    concat_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(235) & concat_CP_34_elements(238);
      gj_concat_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: 	298 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Update/cr
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_update_start_
      -- 
    cr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(237), ack => type_cast_610_inst_req_1); -- 
    concat_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(239) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	233 
    -- CP-element group 238: 	236 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Sample/ra
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_sample_completed_
      -- 
    ra_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_0, ack => concat_CP_34_elements(238)); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	296 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Update/ca
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_610_update_completed_
      -- 
    ca_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_1, ack => concat_CP_34_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	235 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	243 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Sample/rr
      -- CP-element group 240: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_sample_start_
      -- 
    rr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(240), ack => RPIPE_Concat_input_pipe_619_inst_req_0); -- 
    concat_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(235) & concat_CP_34_elements(243);
      gj_concat_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	242 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	246 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_update_start_
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Update/cr
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Update/$entry
      -- 
    cr_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(241), ack => RPIPE_Concat_input_pipe_619_inst_req_1); -- 
    concat_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(242) & concat_CP_34_elements(246);
      gj_concat_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	241 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Sample/ra
      -- 
    ra_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_619_inst_ack_0, ack => concat_CP_34_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: 	248 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	240 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_619_Update/ca
      -- 
    ca_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_619_inst_ack_1, ack => concat_CP_34_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Sample/rr
      -- 
    rr_1267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(244), ack => type_cast_623_inst_req_0); -- 
    concat_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(243) & concat_CP_34_elements(246);
      gj_concat_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: 	298 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_update_start_
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Update/cr
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Update/$entry
      -- 
    cr_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(245), ack => type_cast_623_inst_req_1); -- 
    concat_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(247) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	241 
    -- CP-element group 246: 	244 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Sample/ra
      -- 
    ra_1268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_0, ack => concat_CP_34_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	296 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Update/ca
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_623_Update/$exit
      -- 
    ca_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_1, ack => concat_CP_34_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	243 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	251 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Sample/rr
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Sample/$entry
      -- 
    rr_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(248), ack => RPIPE_Concat_input_pipe_637_inst_req_0); -- 
    concat_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(243) & concat_CP_34_elements(251);
      gj_concat_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	250 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	254 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_update_start_
      -- 
    cr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(249), ack => RPIPE_Concat_input_pipe_637_inst_req_1); -- 
    concat_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(250) & concat_CP_34_elements(254);
      gj_concat_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	249 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Sample/ra
      -- CP-element group 250: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Sample/$exit
      -- 
    ra_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_637_inst_ack_0, ack => concat_CP_34_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251: 	256 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	248 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_Update/ca
      -- CP-element group 251: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_637_update_completed_
      -- 
    ca_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_637_inst_ack_1, ack => concat_CP_34_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Sample/rr
      -- CP-element group 252: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_sample_start_
      -- 
    rr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(252), ack => type_cast_641_inst_req_0); -- 
    concat_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(251) & concat_CP_34_elements(254);
      gj_concat_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	298 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_update_start_
      -- CP-element group 253: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Update/cr
      -- CP-element group 253: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Update/$entry
      -- 
    cr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(253), ack => type_cast_641_inst_req_1); -- 
    concat_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(255) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	249 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Sample/ra
      -- 
    ra_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_0, ack => concat_CP_34_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	296 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Update/ca
      -- CP-element group 255: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_641_Update/$exit
      -- 
    ca_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_1, ack => concat_CP_34_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	251 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	259 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Sample/rr
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_sample_start_
      -- 
    rr_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(256), ack => RPIPE_Concat_input_pipe_655_inst_req_0); -- 
    concat_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(251) & concat_CP_34_elements(259);
      gj_concat_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	258 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	262 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_update_start_
      -- CP-element group 257: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Update/cr
      -- CP-element group 257: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Update/$entry
      -- 
    cr_1314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(257), ack => RPIPE_Concat_input_pipe_655_inst_req_1); -- 
    concat_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(258) & concat_CP_34_elements(262);
      gj_concat_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	257 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Sample/ra
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_sample_completed_
      -- 
    ra_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_655_inst_ack_0, ack => concat_CP_34_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259: 	264 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	256 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_655_update_completed_
      -- 
    ca_1315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_655_inst_ack_1, ack => concat_CP_34_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Sample/rr
      -- 
    rr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(260), ack => type_cast_659_inst_req_0); -- 
    concat_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(259) & concat_CP_34_elements(262);
      gj_concat_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: 	298 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_update_start_
      -- CP-element group 261: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Update/cr
      -- 
    cr_1328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(261), ack => type_cast_659_inst_req_1); -- 
    concat_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(263) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Sample/ra
      -- 
    ra_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_0, ack => concat_CP_34_elements(262)); -- 
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	296 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_659_Update/ca
      -- 
    ca_1329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_1, ack => concat_CP_34_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	259 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	267 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Sample/rr
      -- 
    rr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(264), ack => RPIPE_Concat_input_pipe_673_inst_req_0); -- 
    concat_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(259) & concat_CP_34_elements(267);
      gj_concat_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	266 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	270 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_update_start_
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Update/cr
      -- 
    cr_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(265), ack => RPIPE_Concat_input_pipe_673_inst_req_1); -- 
    concat_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(266) & concat_CP_34_elements(270);
      gj_concat_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	265 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Sample/ra
      -- 
    ra_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_673_inst_ack_0, ack => concat_CP_34_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267: 	272 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	264 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_673_Update/ca
      -- 
    ca_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_673_inst_ack_1, ack => concat_CP_34_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Sample/rr
      -- 
    rr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(268), ack => type_cast_677_inst_req_0); -- 
    concat_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(267) & concat_CP_34_elements(270);
      gj_concat_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	298 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_update_start_
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Update/cr
      -- 
    cr_1356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(269), ack => type_cast_677_inst_req_1); -- 
    concat_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(271) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	265 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Sample/ra
      -- 
    ra_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_0, ack => concat_CP_34_elements(270)); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	296 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_677_Update/ca
      -- 
    ca_1357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_1, ack => concat_CP_34_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	267 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	275 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Sample/rr
      -- 
    rr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(272), ack => RPIPE_Concat_input_pipe_691_inst_req_0); -- 
    concat_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(267) & concat_CP_34_elements(275);
      gj_concat_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	274 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	278 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_update_start_
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Update/cr
      -- 
    cr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(273), ack => RPIPE_Concat_input_pipe_691_inst_req_1); -- 
    concat_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(274) & concat_CP_34_elements(278);
      gj_concat_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	273 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Sample/ra
      -- 
    ra_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_691_inst_ack_0, ack => concat_CP_34_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275: 	280 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	272 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_691_Update/ca
      -- 
    ca_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_691_inst_ack_1, ack => concat_CP_34_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Sample/rr
      -- 
    rr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(276), ack => type_cast_695_inst_req_0); -- 
    concat_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(275) & concat_CP_34_elements(278);
      gj_concat_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: 	298 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_update_start_
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Update/cr
      -- 
    cr_1384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(277), ack => type_cast_695_inst_req_1); -- 
    concat_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(279) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	273 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Sample/ra
      -- 
    ra_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_0, ack => concat_CP_34_elements(278)); -- 
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	296 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_695_Update/ca
      -- 
    ca_1385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_1, ack => concat_CP_34_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	275 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	283 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Sample/rr
      -- 
    rr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(280), ack => RPIPE_Concat_input_pipe_709_inst_req_0); -- 
    concat_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(275) & concat_CP_34_elements(283);
      gj_concat_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	282 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	286 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_update_start_
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Update/cr
      -- 
    cr_1398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(281), ack => RPIPE_Concat_input_pipe_709_inst_req_1); -- 
    concat_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(282) & concat_CP_34_elements(286);
      gj_concat_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	281 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_sample_completed_
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Sample/ra
      -- 
    ra_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_709_inst_ack_0, ack => concat_CP_34_elements(282)); -- 
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283: 	288 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	280 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_709_Update/ca
      -- 
    ca_1399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_709_inst_ack_1, ack => concat_CP_34_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Sample/rr
      -- 
    rr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(284), ack => type_cast_713_inst_req_0); -- 
    concat_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(283) & concat_CP_34_elements(286);
      gj_concat_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: 	298 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_update_start_
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Update/cr
      -- 
    cr_1412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(285), ack => type_cast_713_inst_req_1); -- 
    concat_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(287) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	281 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Sample/ra
      -- 
    ra_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_713_inst_ack_0, ack => concat_CP_34_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	296 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_713_Update/ca
      -- 
    ca_1413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_713_inst_ack_1, ack => concat_CP_34_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	283 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	291 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Sample/rr
      -- 
    rr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(288), ack => RPIPE_Concat_input_pipe_727_inst_req_0); -- 
    concat_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(283) & concat_CP_34_elements(291);
      gj_concat_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	290 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	294 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_update_start_
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Update/cr
      -- 
    cr_1426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(289), ack => RPIPE_Concat_input_pipe_727_inst_req_1); -- 
    concat_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(290) & concat_CP_34_elements(294);
      gj_concat_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	289 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Sample/ra
      -- 
    ra_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_727_inst_ack_0, ack => concat_CP_34_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	233 
    -- CP-element group 291: 	288 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/RPIPE_Concat_input_pipe_727_Update/ca
      -- 
    ca_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_727_inst_ack_1, ack => concat_CP_34_elements(291)); -- 
    -- CP-element group 292:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: marked-predecessors 
    -- CP-element group 292: 	294 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Sample/rr
      -- 
    rr_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(292), ack => type_cast_731_inst_req_0); -- 
    concat_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(291) & concat_CP_34_elements(294);
      gj_concat_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: 	298 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_update_start_
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Update/cr
      -- 
    cr_1440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(293), ack => type_cast_731_inst_req_1); -- 
    concat_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(295) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: successors 
    -- CP-element group 294: marked-successors 
    -- CP-element group 294: 	289 
    -- CP-element group 294: 	292 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_sample_completed_
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Sample/ra
      -- 
    ra_1436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_0, ack => concat_CP_34_elements(294)); -- 
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_update_completed_
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/type_cast_731_Update/ca
      -- 
    ca_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_1, ack => concat_CP_34_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	231 
    -- CP-element group 296: 	239 
    -- CP-element group 296: 	247 
    -- CP-element group 296: 	255 
    -- CP-element group 296: 	263 
    -- CP-element group 296: 	271 
    -- CP-element group 296: 	279 
    -- CP-element group 296: 	287 
    -- CP-element group 296: 	295 
    -- CP-element group 296: marked-predecessors 
    -- CP-element group 296: 	298 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (9) 
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/ptr_deref_739_Split/$entry
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/ptr_deref_739_Split/$exit
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/ptr_deref_739_Split/split_req
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/ptr_deref_739_Split/split_ack
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/word_access_start/$entry
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/word_access_start/word_0/$entry
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/word_access_start/word_0/rr
      -- 
    rr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(296), ack => ptr_deref_739_store_0_req_0); -- 
    concat_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= concat_CP_34_elements(231) & concat_CP_34_elements(239) & concat_CP_34_elements(247) & concat_CP_34_elements(255) & concat_CP_34_elements(263) & concat_CP_34_elements(271) & concat_CP_34_elements(279) & concat_CP_34_elements(287) & concat_CP_34_elements(295) & concat_CP_34_elements(298);
      gj_concat_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (5) 
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_update_start_
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/word_access_complete/$entry
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/word_access_complete/word_0/$entry
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/word_access_complete/word_0/cr
      -- 
    cr_1490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(297), ack => ptr_deref_739_store_0_req_1); -- 
    concat_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(299);
      gj_concat_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: successors 
    -- CP-element group 298: marked-successors 
    -- CP-element group 298: 	226 
    -- CP-element group 298: 	237 
    -- CP-element group 298: 	245 
    -- CP-element group 298: 	253 
    -- CP-element group 298: 	261 
    -- CP-element group 298: 	269 
    -- CP-element group 298: 	277 
    -- CP-element group 298: 	285 
    -- CP-element group 298: 	293 
    -- CP-element group 298: 	296 
    -- CP-element group 298:  members (5) 
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_sample_completed_
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/$exit
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/word_access_start/$exit
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/word_access_start/word_0/$exit
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Sample/word_access_start/word_0/ra
      -- 
    ra_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_739_store_0_ack_0, ack => concat_CP_34_elements(298)); -- 
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (5) 
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_update_completed_
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/$exit
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/word_access_complete/$exit
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/word_access_complete/word_0/$exit
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/ptr_deref_739_Update/word_access_complete/word_0/ca
      -- 
    ca_1491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_739_store_0_ack_1, ack => concat_CP_34_elements(299)); -- 
    -- CP-element group 300:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	203 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	204 
    -- CP-element group 300:  members (1) 
      -- CP-element group 300: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group concat_CP_34_elements(300) is a control-delay.
    cp_element_300_delay: control_delay_element  generic map(name => " 300_delay", delay_value => 1)  port map(req => concat_CP_34_elements(203), ack => concat_CP_34_elements(300), clk => clk, reset =>reset);
    -- CP-element group 301:  join  transition  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	208 
    -- CP-element group 301: 	228 
    -- CP-element group 301: 	299 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	200 
    -- CP-element group 301:  members (1) 
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_590/do_while_stmt_590_loop_body/$exit
      -- 
    concat_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(208) & concat_CP_34_elements(228) & concat_CP_34_elements(299);
      gj_concat_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	199 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (2) 
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_590/loop_exit/$exit
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_590/loop_exit/ack
      -- 
    ack_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_590_branch_ack_0, ack => concat_CP_34_elements(302)); -- 
    -- CP-element group 303:  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	199 
    -- CP-element group 303: successors 
    -- CP-element group 303:  members (2) 
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_590/loop_taken/$exit
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_590/loop_taken/ack
      -- 
    ack_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_590_branch_ack_1, ack => concat_CP_34_elements(303)); -- 
    -- CP-element group 304:  transition  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	197 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	2 
    -- CP-element group 304:  members (1) 
      -- CP-element group 304: 	 branch_block_stmt_23/do_while_stmt_590/$exit
      -- 
    concat_CP_34_elements(304) <= concat_CP_34_elements(197);
    -- CP-element group 305:  merge  transition  place  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	2 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	795 
    -- CP-element group 305:  members (13) 
      -- CP-element group 305: 	 branch_block_stmt_23/merge_stmt_763__exit__
      -- CP-element group 305: 	 branch_block_stmt_23/forx_xend223x_xloopexit_forx_xend223
      -- CP-element group 305: 	 branch_block_stmt_23/if_stmt_759_if_link/$exit
      -- CP-element group 305: 	 branch_block_stmt_23/if_stmt_759_if_link/if_choice_transition
      -- CP-element group 305: 	 branch_block_stmt_23/forx_xbody169_forx_xend223x_xloopexit
      -- CP-element group 305: 	 branch_block_stmt_23/forx_xbody169_forx_xend223x_xloopexit_PhiReq/$entry
      -- CP-element group 305: 	 branch_block_stmt_23/forx_xbody169_forx_xend223x_xloopexit_PhiReq/$exit
      -- CP-element group 305: 	 branch_block_stmt_23/merge_stmt_763_PhiReqMerge
      -- CP-element group 305: 	 branch_block_stmt_23/merge_stmt_763_PhiAck/$entry
      -- CP-element group 305: 	 branch_block_stmt_23/merge_stmt_763_PhiAck/$exit
      -- CP-element group 305: 	 branch_block_stmt_23/merge_stmt_763_PhiAck/dummy
      -- CP-element group 305: 	 branch_block_stmt_23/forx_xend223x_xloopexit_forx_xend223_PhiReq/$entry
      -- CP-element group 305: 	 branch_block_stmt_23/forx_xend223x_xloopexit_forx_xend223_PhiReq/$exit
      -- 
    if_choice_transition_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_759_branch_ack_1, ack => concat_CP_34_elements(305)); -- 
    -- CP-element group 306:  merge  transition  place  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	2 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (5) 
      -- CP-element group 306: 	 branch_block_stmt_23/if_stmt_759__exit__
      -- CP-element group 306: 	 branch_block_stmt_23/merge_stmt_763__entry__
      -- CP-element group 306: 	 branch_block_stmt_23/if_stmt_759_else_link/$exit
      -- CP-element group 306: 	 branch_block_stmt_23/if_stmt_759_else_link/else_choice_transition
      -- CP-element group 306: 	 branch_block_stmt_23/merge_stmt_763_dead_link/$entry
      -- 
    else_choice_transition_1518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_759_branch_ack_0, ack => concat_CP_34_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	795 
    -- CP-element group 307: successors 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/cra
      -- 
    cra_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_768_call_ack_0, ack => concat_CP_34_elements(307)); -- 
    -- CP-element group 308:  transition  place  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	795 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (17) 
      -- CP-element group 308: 	 branch_block_stmt_23/call_stmt_768__exit__
      -- CP-element group 308: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787__entry__
      -- CP-element group 308: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787__exit__
      -- CP-element group 308: 	 branch_block_stmt_23/forx_xend223_whilex_xbody
      -- CP-element group 308: 	 branch_block_stmt_23/merge_stmt_789__exit__
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_817__entry__
      -- CP-element group 308: 	 branch_block_stmt_23/call_stmt_768/$exit
      -- CP-element group 308: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/cca
      -- CP-element group 308: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787/$exit
      -- CP-element group 308: 	 branch_block_stmt_23/forx_xend223_whilex_xbody_PhiReq/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/forx_xend223_whilex_xbody_PhiReq/$exit
      -- CP-element group 308: 	 branch_block_stmt_23/merge_stmt_789_PhiReqMerge
      -- CP-element group 308: 	 branch_block_stmt_23/merge_stmt_789_PhiAck/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/merge_stmt_789_PhiAck/$exit
      -- 
    cca_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_768_call_ack_1, ack => concat_CP_34_elements(308)); -- 
    -- CP-element group 309:  transition  place  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	315 
    -- CP-element group 309:  members (2) 
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_817/$entry
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817__entry__
      -- 
    concat_CP_34_elements(309) <= concat_CP_34_elements(308);
    -- CP-element group 310:  merge  place  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	694 
    -- CP-element group 310:  members (1) 
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817__exit__
      -- 
    -- Element group concat_CP_34_elements(310) is bound as output of CP function.
    -- CP-element group 311:  merge  place  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	314 
    -- CP-element group 311:  members (1) 
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/loop_back
      -- 
    -- Element group concat_CP_34_elements(311) is bound as output of CP function.
    -- CP-element group 312:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	317 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	692 
    -- CP-element group 312: 	693 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_817/condition_done
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_817/loop_exit/$entry
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_817/loop_taken/$entry
      -- 
    concat_CP_34_elements(312) <= concat_CP_34_elements(317);
    -- CP-element group 313:  branch  place  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	691 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_23/do_while_stmt_817/loop_body_done
      -- 
    concat_CP_34_elements(313) <= concat_CP_34_elements(691);
    -- CP-element group 314:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	311 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	347 
    -- CP-element group 314: 	368 
    -- CP-element group 314: 	389 
    -- CP-element group 314: 	410 
    -- CP-element group 314: 	328 
    -- CP-element group 314:  members (1) 
      -- CP-element group 314: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/back_edge_to_loop_body
      -- 
    concat_CP_34_elements(314) <= concat_CP_34_elements(311);
    -- CP-element group 315:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	309 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	349 
    -- CP-element group 315: 	370 
    -- CP-element group 315: 	391 
    -- CP-element group 315: 	412 
    -- CP-element group 315: 	330 
    -- CP-element group 315:  members (1) 
      -- CP-element group 315: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/first_time_through_loop_body
      -- 
    concat_CP_34_elements(315) <= concat_CP_34_elements(309);
    -- CP-element group 316:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	343 
    -- CP-element group 316: 	344 
    -- CP-element group 316: 	362 
    -- CP-element group 316: 	363 
    -- CP-element group 316: 	383 
    -- CP-element group 316: 	384 
    -- CP-element group 316: 	404 
    -- CP-element group 316: 	405 
    -- CP-element group 316: 	438 
    -- CP-element group 316: 	439 
    -- CP-element group 316: 	461 
    -- CP-element group 316: 	462 
    -- CP-element group 316: 	548 
    -- CP-element group 316: 	549 
    -- CP-element group 316: 	571 
    -- CP-element group 316: 	572 
    -- CP-element group 316: 	689 
    -- CP-element group 316: 	322 
    -- CP-element group 316: 	323 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/$entry
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/loop_body_start
      -- 
    -- Element group concat_CP_34_elements(316) is bound as output of CP function.
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	688 
    -- CP-element group 317: 	689 
    -- CP-element group 317: 	321 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	312 
    -- CP-element group 317:  members (1) 
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/condition_evaluated
      -- 
    condition_evaluated_1554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(317), ack => do_while_stmt_817_branch_req_0); -- 
    concat_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(688) & concat_CP_34_elements(689) & concat_CP_34_elements(321);
      gj_concat_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	343 
    -- CP-element group 318: 	362 
    -- CP-element group 318: 	383 
    -- CP-element group 318: 	404 
    -- CP-element group 318: 	322 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	321 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	364 
    -- CP-element group 318: 	385 
    -- CP-element group 318: 	406 
    -- CP-element group 318: 	324 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_sample_req
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_start__ps
      -- 
    concat_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(343) & concat_CP_34_elements(362) & concat_CP_34_elements(383) & concat_CP_34_elements(404) & concat_CP_34_elements(322) & concat_CP_34_elements(321);
      gj_concat_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	345 
    -- CP-element group 319: 	365 
    -- CP-element group 319: 	386 
    -- CP-element group 319: 	407 
    -- CP-element group 319: 	325 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	426 
    -- CP-element group 319: 	484 
    -- CP-element group 319: 	496 
    -- CP-element group 319: 	614 
    -- CP-element group 319: 	622 
    -- CP-element group 319: 	626 
    -- CP-element group 319: 	630 
    -- CP-element group 319: 	634 
    -- CP-element group 319: 	642 
    -- CP-element group 319: 	646 
    -- CP-element group 319: 	650 
    -- CP-element group 319: 	658 
    -- CP-element group 319: 	662 
    -- CP-element group 319: 	670 
    -- CP-element group 319: 	674 
    -- CP-element group 319: 	682 
    -- CP-element group 319: marked-successors 
    -- CP-element group 319: 	343 
    -- CP-element group 319: 	362 
    -- CP-element group 319: 	383 
    -- CP-element group 319: 	404 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (6) 
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_sample_ack
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_completed_
      -- 
    concat_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(345) & concat_CP_34_elements(365) & concat_CP_34_elements(386) & concat_CP_34_elements(407) & concat_CP_34_elements(325);
      gj_concat_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	344 
    -- CP-element group 320: 	363 
    -- CP-element group 320: 	384 
    -- CP-element group 320: 	405 
    -- CP-element group 320: 	323 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	366 
    -- CP-element group 320: 	387 
    -- CP-element group 320: 	408 
    -- CP-element group 320: 	326 
    -- CP-element group 320:  members (2) 
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_update_req
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_start__ps
      -- 
    concat_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(344) & concat_CP_34_elements(363) & concat_CP_34_elements(384) & concat_CP_34_elements(405) & concat_CP_34_elements(323);
      gj_concat_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	346 
    -- CP-element group 321: 	367 
    -- CP-element group 321: 	388 
    -- CP-element group 321: 	409 
    -- CP-element group 321: 	327 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	317 
    -- CP-element group 321: marked-successors 
    -- CP-element group 321: 	318 
    -- CP-element group 321:  members (1) 
      -- CP-element group 321: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_update_ack
      -- 
    concat_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(346) & concat_CP_34_elements(367) & concat_CP_34_elements(388) & concat_CP_34_elements(409) & concat_CP_34_elements(327);
      gj_concat_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	316 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	616 
    -- CP-element group 322: 	624 
    -- CP-element group 322: 	628 
    -- CP-element group 322: 	648 
    -- CP-element group 322: 	652 
    -- CP-element group 322: 	660 
    -- CP-element group 322: 	319 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	318 
    -- CP-element group 322:  members (1) 
      -- CP-element group 322: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_start_
      -- 
    concat_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(616) & concat_CP_34_elements(624) & concat_CP_34_elements(628) & concat_CP_34_elements(648) & concat_CP_34_elements(652) & concat_CP_34_elements(660) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  join  transition  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	316 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	454 
    -- CP-element group 323: 	489 
    -- CP-element group 323: 	493 
    -- CP-element group 323: 	327 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	320 
    -- CP-element group 323:  members (1) 
      -- CP-element group 323: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_start_
      -- 
    concat_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(454) & concat_CP_34_elements(489) & concat_CP_34_elements(493) & concat_CP_34_elements(327);
      gj_concat_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	318 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (1) 
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_start__ps
      -- 
    concat_CP_34_elements(324) <= concat_CP_34_elements(318);
    -- CP-element group 325:  join  transition  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	319 
    -- CP-element group 325:  members (1) 
      -- CP-element group 325: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(325) is bound as output of CP function.
    -- CP-element group 326:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	320 
    -- CP-element group 326: successors 
    -- CP-element group 326:  members (1) 
      -- CP-element group 326: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_start__ps
      -- 
    concat_CP_34_elements(326) <= concat_CP_34_elements(320);
    -- CP-element group 327:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	452 
    -- CP-element group 327: 	487 
    -- CP-element group 327: 	491 
    -- CP-element group 327: 	321 
    -- CP-element group 327: marked-successors 
    -- CP-element group 327: 	323 
    -- CP-element group 327:  members (2) 
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_completed_
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(327) is bound as output of CP function.
    -- CP-element group 328:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	314 
    -- CP-element group 328: successors 
    -- CP-element group 328:  members (1) 
      -- CP-element group 328: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_loopback_trigger
      -- 
    concat_CP_34_elements(328) <= concat_CP_34_elements(314);
    -- CP-element group 329:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: successors 
    -- CP-element group 329:  members (2) 
      -- CP-element group 329: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_loopback_sample_req
      -- CP-element group 329: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_loopback_sample_req_ps
      -- 
    phi_stmt_819_loopback_sample_req_1569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_819_loopback_sample_req_1569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(329), ack => phi_stmt_819_req_0); -- 
    -- Element group concat_CP_34_elements(329) is bound as output of CP function.
    -- CP-element group 330:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	315 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_entry_trigger
      -- 
    concat_CP_34_elements(330) <= concat_CP_34_elements(315);
    -- CP-element group 331:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: successors 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_entry_sample_req
      -- CP-element group 331: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_entry_sample_req_ps
      -- 
    phi_stmt_819_entry_sample_req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_819_entry_sample_req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(331), ack => phi_stmt_819_req_1); -- 
    -- Element group concat_CP_34_elements(331) is bound as output of CP function.
    -- CP-element group 332:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_phi_mux_ack
      -- CP-element group 332: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_phi_mux_ack_ps
      -- 
    phi_stmt_819_phi_mux_ack_1575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_819_ack_0, ack => concat_CP_34_elements(332)); -- 
    -- CP-element group 333:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (1) 
      -- CP-element group 333: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(333) is bound as output of CP function.
    -- CP-element group 334:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (1) 
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(334) is bound as output of CP function.
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/rr
      -- 
    rr_1588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(335), ack => type_cast_822_inst_req_0); -- 
    concat_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(333) & concat_CP_34_elements(337);
      gj_concat_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: marked-predecessors 
    -- CP-element group 336: 	338 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	338 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_start_
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/cr
      -- 
    cr_1593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(336), ack => type_cast_822_inst_req_1); -- 
    concat_cp_element_group_336: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_336"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(334) & concat_CP_34_elements(338);
      gj_concat_cp_element_group_336 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(336), clk => clk, reset => reset); --
    end block;
    -- CP-element group 337:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: marked-successors 
    -- CP-element group 337: 	335 
    -- CP-element group 337:  members (4) 
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_completed__ps
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/ra
      -- 
    ra_1589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_0, ack => concat_CP_34_elements(337)); -- 
    -- CP-element group 338:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: marked-successors 
    -- CP-element group 338: 	336 
    -- CP-element group 338:  members (4) 
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_completed__ps
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/ca
      -- 
    ca_1594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_1, ack => concat_CP_34_elements(338)); -- 
    -- CP-element group 339:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: successors 
    -- CP-element group 339:  members (4) 
      -- CP-element group 339: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_start__ps
      -- CP-element group 339: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_completed__ps
      -- CP-element group 339: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(339) is bound as output of CP function.
    -- CP-element group 340:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (2) 
      -- CP-element group 340: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_start__ps
      -- CP-element group 340: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_start_
      -- 
    -- Element group concat_CP_34_elements(340) is bound as output of CP function.
    -- CP-element group 341:  join  transition  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: successors 
    -- CP-element group 341:  members (1) 
      -- CP-element group 341: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_completed__ps
      -- 
    concat_CP_34_elements(341) <= concat_CP_34_elements(342);
    -- CP-element group 342:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	341 
    -- CP-element group 342:  members (1) 
      -- CP-element group 342: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_completed_
      -- 
    -- Element group concat_CP_34_elements(342) is a control-delay.
    cp_element_342_delay: control_delay_element  generic map(name => " 342_delay", delay_value => 1)  port map(req => concat_CP_34_elements(340), ack => concat_CP_34_elements(342), clk => clk, reset =>reset);
    -- CP-element group 343:  join  transition  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	316 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	428 
    -- CP-element group 343: 	486 
    -- CP-element group 343: 	498 
    -- CP-element group 343: 	319 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	318 
    -- CP-element group 343:  members (1) 
      -- CP-element group 343: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_start_
      -- 
    concat_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(428) & concat_CP_34_elements(486) & concat_CP_34_elements(498) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  join  transition  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	316 
    -- CP-element group 344: marked-predecessors 
    -- CP-element group 344: 	346 
    -- CP-element group 344: 	431 
    -- CP-element group 344: 	485 
    -- CP-element group 344: 	497 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	320 
    -- CP-element group 344:  members (1) 
      -- CP-element group 344: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_start_
      -- 
    concat_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(346) & concat_CP_34_elements(431) & concat_CP_34_elements(485) & concat_CP_34_elements(497);
      gj_concat_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  join  transition  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	319 
    -- CP-element group 345:  members (1) 
      -- CP-element group 345: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(345) is bound as output of CP function.
    -- CP-element group 346:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	429 
    -- CP-element group 346: 	483 
    -- CP-element group 346: 	495 
    -- CP-element group 346: 	321 
    -- CP-element group 346: marked-successors 
    -- CP-element group 346: 	344 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(346) is bound as output of CP function.
    -- CP-element group 347:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	314 
    -- CP-element group 347: successors 
    -- CP-element group 347:  members (1) 
      -- CP-element group 347: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_loopback_trigger
      -- 
    concat_CP_34_elements(347) <= concat_CP_34_elements(314);
    -- CP-element group 348:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (2) 
      -- CP-element group 348: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_loopback_sample_req
      -- CP-element group 348: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_loopback_sample_req_ps
      -- 
    phi_stmt_824_loopback_sample_req_1613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_824_loopback_sample_req_1613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(348), ack => phi_stmt_824_req_0); -- 
    -- Element group concat_CP_34_elements(348) is bound as output of CP function.
    -- CP-element group 349:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	315 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (1) 
      -- CP-element group 349: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_entry_trigger
      -- 
    concat_CP_34_elements(349) <= concat_CP_34_elements(315);
    -- CP-element group 350:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (2) 
      -- CP-element group 350: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_entry_sample_req
      -- CP-element group 350: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_entry_sample_req_ps
      -- 
    phi_stmt_824_entry_sample_req_1616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_824_entry_sample_req_1616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(350), ack => phi_stmt_824_req_1); -- 
    -- Element group concat_CP_34_elements(350) is bound as output of CP function.
    -- CP-element group 351:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: successors 
    -- CP-element group 351:  members (2) 
      -- CP-element group 351: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_phi_mux_ack
      -- CP-element group 351: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_phi_mux_ack_ps
      -- 
    phi_stmt_824_phi_mux_ack_1619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_824_ack_0, ack => concat_CP_34_elements(351)); -- 
    -- CP-element group 352:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	354 
    -- CP-element group 352:  members (1) 
      -- CP-element group 352: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(352) is bound as output of CP function.
    -- CP-element group 353:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (1) 
      -- CP-element group 353: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(353) is bound as output of CP function.
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	352 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/rr
      -- 
    rr_1632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(354), ack => type_cast_827_inst_req_0); -- 
    concat_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(352) & concat_CP_34_elements(356);
      gj_concat_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	357 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_start_
      -- CP-element group 355: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/cr
      -- 
    cr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(355), ack => type_cast_827_inst_req_1); -- 
    concat_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(353) & concat_CP_34_elements(357);
      gj_concat_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (4) 
      -- CP-element group 356: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_completed__ps
      -- CP-element group 356: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/ra
      -- 
    ra_1633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_0, ack => concat_CP_34_elements(356)); -- 
    -- CP-element group 357:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: marked-successors 
    -- CP-element group 357: 	355 
    -- CP-element group 357:  members (4) 
      -- CP-element group 357: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_completed__ps
      -- CP-element group 357: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/ca
      -- 
    ca_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_1, ack => concat_CP_34_elements(357)); -- 
    -- CP-element group 358:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: successors 
    -- CP-element group 358:  members (4) 
      -- CP-element group 358: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_start__ps
      -- CP-element group 358: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_completed__ps
      -- CP-element group 358: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(358) is bound as output of CP function.
    -- CP-element group 359:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (2) 
      -- CP-element group 359: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_start__ps
      -- CP-element group 359: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_start_
      -- 
    -- Element group concat_CP_34_elements(359) is bound as output of CP function.
    -- CP-element group 360:  join  transition  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	361 
    -- CP-element group 360: successors 
    -- CP-element group 360:  members (1) 
      -- CP-element group 360: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_completed__ps
      -- 
    concat_CP_34_elements(360) <= concat_CP_34_elements(361);
    -- CP-element group 361:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	360 
    -- CP-element group 361:  members (1) 
      -- CP-element group 361: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_completed_
      -- 
    -- Element group concat_CP_34_elements(361) is a control-delay.
    cp_element_361_delay: control_delay_element  generic map(name => " 361_delay", delay_value => 1)  port map(req => concat_CP_34_elements(359), ack => concat_CP_34_elements(361), clk => clk, reset =>reset);
    -- CP-element group 362:  join  transition  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	316 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	616 
    -- CP-element group 362: 	624 
    -- CP-element group 362: 	628 
    -- CP-element group 362: 	632 
    -- CP-element group 362: 	636 
    -- CP-element group 362: 	644 
    -- CP-element group 362: 	319 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	318 
    -- CP-element group 362:  members (1) 
      -- CP-element group 362: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_start_
      -- 
    concat_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(616) & concat_CP_34_elements(624) & concat_CP_34_elements(628) & concat_CP_34_elements(632) & concat_CP_34_elements(636) & concat_CP_34_elements(644) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  join  transition  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	316 
    -- CP-element group 363: marked-predecessors 
    -- CP-element group 363: 	367 
    -- CP-element group 363: 	541 
    -- CP-element group 363: 	595 
    -- CP-element group 363: 	607 
    -- CP-element group 363: 	639 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	320 
    -- CP-element group 363:  members (1) 
      -- CP-element group 363: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_start_
      -- 
    concat_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(367) & concat_CP_34_elements(541) & concat_CP_34_elements(595) & concat_CP_34_elements(607) & concat_CP_34_elements(639);
      gj_concat_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	318 
    -- CP-element group 364: successors 
    -- CP-element group 364:  members (1) 
      -- CP-element group 364: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_start__ps
      -- 
    concat_CP_34_elements(364) <= concat_CP_34_elements(318);
    -- CP-element group 365:  join  transition  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	319 
    -- CP-element group 365:  members (1) 
      -- CP-element group 365: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(365) is bound as output of CP function.
    -- CP-element group 366:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	320 
    -- CP-element group 366: successors 
    -- CP-element group 366:  members (1) 
      -- CP-element group 366: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_start__ps
      -- 
    concat_CP_34_elements(366) <= concat_CP_34_elements(320);
    -- CP-element group 367:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	539 
    -- CP-element group 367: 	593 
    -- CP-element group 367: 	605 
    -- CP-element group 367: 	637 
    -- CP-element group 367: 	321 
    -- CP-element group 367: marked-successors 
    -- CP-element group 367: 	363 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(367) is bound as output of CP function.
    -- CP-element group 368:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	314 
    -- CP-element group 368: successors 
    -- CP-element group 368:  members (1) 
      -- CP-element group 368: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_loopback_trigger
      -- 
    concat_CP_34_elements(368) <= concat_CP_34_elements(314);
    -- CP-element group 369:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: successors 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_loopback_sample_req
      -- CP-element group 369: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_loopback_sample_req_ps
      -- 
    phi_stmt_829_loopback_sample_req_1657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_829_loopback_sample_req_1657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(369), ack => phi_stmt_829_req_0); -- 
    -- Element group concat_CP_34_elements(369) is bound as output of CP function.
    -- CP-element group 370:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	315 
    -- CP-element group 370: successors 
    -- CP-element group 370:  members (1) 
      -- CP-element group 370: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_entry_trigger
      -- 
    concat_CP_34_elements(370) <= concat_CP_34_elements(315);
    -- CP-element group 371:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: successors 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_entry_sample_req
      -- CP-element group 371: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_entry_sample_req_ps
      -- 
    phi_stmt_829_entry_sample_req_1660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_829_entry_sample_req_1660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(371), ack => phi_stmt_829_req_1); -- 
    -- Element group concat_CP_34_elements(371) is bound as output of CP function.
    -- CP-element group 372:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: successors 
    -- CP-element group 372:  members (2) 
      -- CP-element group 372: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_phi_mux_ack
      -- CP-element group 372: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_phi_mux_ack_ps
      -- 
    phi_stmt_829_phi_mux_ack_1663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_829_ack_0, ack => concat_CP_34_elements(372)); -- 
    -- CP-element group 373:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (1) 
      -- CP-element group 373: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(373) is bound as output of CP function.
    -- CP-element group 374:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (1) 
      -- CP-element group 374: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(374) is bound as output of CP function.
    -- CP-element group 375:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: marked-predecessors 
    -- CP-element group 375: 	377 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/rr
      -- 
    rr_1676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(375), ack => type_cast_832_inst_req_0); -- 
    concat_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(373) & concat_CP_34_elements(377);
      gj_concat_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_start_
      -- CP-element group 376: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/cr
      -- 
    cr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(376), ack => type_cast_832_inst_req_1); -- 
    concat_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(374) & concat_CP_34_elements(378);
      gj_concat_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: marked-successors 
    -- CP-element group 377: 	375 
    -- CP-element group 377:  members (4) 
      -- CP-element group 377: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_completed__ps
      -- CP-element group 377: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/ra
      -- 
    ra_1677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_0, ack => concat_CP_34_elements(377)); -- 
    -- CP-element group 378:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (4) 
      -- CP-element group 378: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_completed__ps
      -- CP-element group 378: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/ca
      -- 
    ca_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_1, ack => concat_CP_34_elements(378)); -- 
    -- CP-element group 379:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: successors 
    -- CP-element group 379:  members (4) 
      -- CP-element group 379: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_start__ps
      -- CP-element group 379: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_completed__ps
      -- CP-element group 379: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(379) is bound as output of CP function.
    -- CP-element group 380:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (2) 
      -- CP-element group 380: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_start__ps
      -- CP-element group 380: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_start_
      -- 
    -- Element group concat_CP_34_elements(380) is bound as output of CP function.
    -- CP-element group 381:  join  transition  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	382 
    -- CP-element group 381: successors 
    -- CP-element group 381:  members (1) 
      -- CP-element group 381: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_completed__ps
      -- 
    concat_CP_34_elements(381) <= concat_CP_34_elements(382);
    -- CP-element group 382:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	381 
    -- CP-element group 382:  members (1) 
      -- CP-element group 382: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_completed_
      -- 
    -- Element group concat_CP_34_elements(382) is a control-delay.
    cp_element_382_delay: control_delay_element  generic map(name => " 382_delay", delay_value => 1)  port map(req => concat_CP_34_elements(380), ack => concat_CP_34_elements(382), clk => clk, reset =>reset);
    -- CP-element group 383:  join  transition  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	316 
    -- CP-element group 383: marked-predecessors 
    -- CP-element group 383: 	616 
    -- CP-element group 383: 	624 
    -- CP-element group 383: 	628 
    -- CP-element group 383: 	664 
    -- CP-element group 383: 	672 
    -- CP-element group 383: 	319 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	318 
    -- CP-element group 383:  members (1) 
      -- CP-element group 383: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_start_
      -- 
    concat_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(616) & concat_CP_34_elements(624) & concat_CP_34_elements(628) & concat_CP_34_elements(664) & concat_CP_34_elements(672) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  join  transition  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	316 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	388 
    -- CP-element group 384: 	427 
    -- CP-element group 384: 	481 
    -- CP-element group 384: 	501 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	320 
    -- CP-element group 384:  members (1) 
      -- CP-element group 384: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_start_
      -- 
    concat_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(388) & concat_CP_34_elements(427) & concat_CP_34_elements(481) & concat_CP_34_elements(501);
      gj_concat_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	318 
    -- CP-element group 385: successors 
    -- CP-element group 385:  members (1) 
      -- CP-element group 385: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_start__ps
      -- 
    concat_CP_34_elements(385) <= concat_CP_34_elements(318);
    -- CP-element group 386:  join  transition  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	319 
    -- CP-element group 386:  members (1) 
      -- CP-element group 386: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(386) is bound as output of CP function.
    -- CP-element group 387:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	320 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (1) 
      -- CP-element group 387: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_start__ps
      -- 
    concat_CP_34_elements(387) <= concat_CP_34_elements(320);
    -- CP-element group 388:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	425 
    -- CP-element group 388: 	479 
    -- CP-element group 388: 	499 
    -- CP-element group 388: 	321 
    -- CP-element group 388: marked-successors 
    -- CP-element group 388: 	384 
    -- CP-element group 388:  members (2) 
      -- CP-element group 388: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(388) is bound as output of CP function.
    -- CP-element group 389:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	314 
    -- CP-element group 389: successors 
    -- CP-element group 389:  members (1) 
      -- CP-element group 389: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_loopback_trigger
      -- 
    concat_CP_34_elements(389) <= concat_CP_34_elements(314);
    -- CP-element group 390:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (2) 
      -- CP-element group 390: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_loopback_sample_req
      -- CP-element group 390: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_loopback_sample_req_ps
      -- 
    phi_stmt_834_loopback_sample_req_1701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_834_loopback_sample_req_1701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(390), ack => phi_stmt_834_req_0); -- 
    -- Element group concat_CP_34_elements(390) is bound as output of CP function.
    -- CP-element group 391:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	315 
    -- CP-element group 391: successors 
    -- CP-element group 391:  members (1) 
      -- CP-element group 391: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_entry_trigger
      -- 
    concat_CP_34_elements(391) <= concat_CP_34_elements(315);
    -- CP-element group 392:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (2) 
      -- CP-element group 392: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_entry_sample_req
      -- CP-element group 392: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_entry_sample_req_ps
      -- 
    phi_stmt_834_entry_sample_req_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_834_entry_sample_req_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(392), ack => phi_stmt_834_req_1); -- 
    -- Element group concat_CP_34_elements(392) is bound as output of CP function.
    -- CP-element group 393:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (2) 
      -- CP-element group 393: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_phi_mux_ack_ps
      -- CP-element group 393: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_phi_mux_ack
      -- 
    phi_stmt_834_phi_mux_ack_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_834_ack_0, ack => concat_CP_34_elements(393)); -- 
    -- CP-element group 394:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	396 
    -- CP-element group 394:  members (1) 
      -- CP-element group 394: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(394) is bound as output of CP function.
    -- CP-element group 395:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(395) is bound as output of CP function.
    -- CP-element group 396:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	394 
    -- CP-element group 396: marked-predecessors 
    -- CP-element group 396: 	398 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	398 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_start_
      -- 
    rr_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_837_inst_req_0); -- 
    concat_cp_element_group_396: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_396"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(394) & concat_CP_34_elements(398);
      gj_concat_cp_element_group_396 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(396), clk => clk, reset => reset); --
    end block;
    -- CP-element group 397:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: marked-predecessors 
    -- CP-element group 397: 	399 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	399 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/cr
      -- CP-element group 397: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_start_
      -- 
    cr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(397), ack => type_cast_837_inst_req_1); -- 
    concat_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(395) & concat_CP_34_elements(399);
      gj_concat_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	396 
    -- CP-element group 398: successors 
    -- CP-element group 398: marked-successors 
    -- CP-element group 398: 	396 
    -- CP-element group 398:  members (4) 
      -- CP-element group 398: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/ra
      -- CP-element group 398: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_completed__ps
      -- 
    ra_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_0, ack => concat_CP_34_elements(398)); -- 
    -- CP-element group 399:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	397 
    -- CP-element group 399: successors 
    -- CP-element group 399: marked-successors 
    -- CP-element group 399: 	397 
    -- CP-element group 399:  members (4) 
      -- CP-element group 399: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/ca
      -- CP-element group 399: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_completed__ps
      -- 
    ca_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_1, ack => concat_CP_34_elements(399)); -- 
    -- CP-element group 400:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: successors 
    -- CP-element group 400:  members (4) 
      -- CP-element group 400: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_start__ps
      -- CP-element group 400: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_completed__ps
      -- CP-element group 400: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(400) is bound as output of CP function.
    -- CP-element group 401:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	403 
    -- CP-element group 401:  members (2) 
      -- CP-element group 401: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_start_
      -- CP-element group 401: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(401) is bound as output of CP function.
    -- CP-element group 402:  join  transition  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	403 
    -- CP-element group 402: successors 
    -- CP-element group 402:  members (1) 
      -- CP-element group 402: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_completed__ps
      -- 
    concat_CP_34_elements(402) <= concat_CP_34_elements(403);
    -- CP-element group 403:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	401 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	402 
    -- CP-element group 403:  members (1) 
      -- CP-element group 403: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_completed_
      -- 
    -- Element group concat_CP_34_elements(403) is a control-delay.
    cp_element_403_delay: control_delay_element  generic map(name => " 403_delay", delay_value => 1)  port map(req => concat_CP_34_elements(401), ack => concat_CP_34_elements(403), clk => clk, reset =>reset);
    -- CP-element group 404:  join  transition  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	316 
    -- CP-element group 404: marked-predecessors 
    -- CP-element group 404: 	616 
    -- CP-element group 404: 	624 
    -- CP-element group 404: 	628 
    -- CP-element group 404: 	676 
    -- CP-element group 404: 	684 
    -- CP-element group 404: 	319 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	318 
    -- CP-element group 404:  members (1) 
      -- CP-element group 404: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_start_
      -- 
    concat_cp_element_group_404: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_404"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(616) & concat_CP_34_elements(624) & concat_CP_34_elements(628) & concat_CP_34_elements(676) & concat_CP_34_elements(684) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_404 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(404), clk => clk, reset => reset); --
    end block;
    -- CP-element group 405:  join  transition  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	316 
    -- CP-element group 405: marked-predecessors 
    -- CP-element group 405: 	409 
    -- CP-element group 405: 	521 
    -- CP-element group 405: 	591 
    -- CP-element group 405: 	611 
    -- CP-element group 405: 	679 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	320 
    -- CP-element group 405:  members (1) 
      -- CP-element group 405: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_start_
      -- 
    concat_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(409) & concat_CP_34_elements(521) & concat_CP_34_elements(591) & concat_CP_34_elements(611) & concat_CP_34_elements(679);
      gj_concat_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	318 
    -- CP-element group 406: successors 
    -- CP-element group 406:  members (1) 
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_start__ps
      -- 
    concat_CP_34_elements(406) <= concat_CP_34_elements(318);
    -- CP-element group 407:  join  transition  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	319 
    -- CP-element group 407:  members (1) 
      -- CP-element group 407: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(407) is bound as output of CP function.
    -- CP-element group 408:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	320 
    -- CP-element group 408: successors 
    -- CP-element group 408:  members (1) 
      -- CP-element group 408: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_start__ps
      -- 
    concat_CP_34_elements(408) <= concat_CP_34_elements(320);
    -- CP-element group 409:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	519 
    -- CP-element group 409: 	589 
    -- CP-element group 409: 	609 
    -- CP-element group 409: 	677 
    -- CP-element group 409: 	321 
    -- CP-element group 409: marked-successors 
    -- CP-element group 409: 	405 
    -- CP-element group 409:  members (2) 
      -- CP-element group 409: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_completed_
      -- CP-element group 409: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(409) is bound as output of CP function.
    -- CP-element group 410:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	314 
    -- CP-element group 410: successors 
    -- CP-element group 410:  members (1) 
      -- CP-element group 410: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_loopback_trigger
      -- 
    concat_CP_34_elements(410) <= concat_CP_34_elements(314);
    -- CP-element group 411:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: successors 
    -- CP-element group 411:  members (2) 
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_loopback_sample_req
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_loopback_sample_req_ps
      -- 
    phi_stmt_839_loopback_sample_req_1745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_839_loopback_sample_req_1745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(411), ack => phi_stmt_839_req_0); -- 
    -- Element group concat_CP_34_elements(411) is bound as output of CP function.
    -- CP-element group 412:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	315 
    -- CP-element group 412: successors 
    -- CP-element group 412:  members (1) 
      -- CP-element group 412: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_entry_trigger
      -- 
    concat_CP_34_elements(412) <= concat_CP_34_elements(315);
    -- CP-element group 413:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: successors 
    -- CP-element group 413:  members (2) 
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_entry_sample_req_ps
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_entry_sample_req
      -- 
    phi_stmt_839_entry_sample_req_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_839_entry_sample_req_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(413), ack => phi_stmt_839_req_1); -- 
    -- Element group concat_CP_34_elements(413) is bound as output of CP function.
    -- CP-element group 414:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: successors 
    -- CP-element group 414:  members (2) 
      -- CP-element group 414: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_phi_mux_ack
      -- CP-element group 414: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_phi_mux_ack_ps
      -- 
    phi_stmt_839_phi_mux_ack_1751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_839_ack_0, ack => concat_CP_34_elements(414)); -- 
    -- CP-element group 415:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	417 
    -- CP-element group 415:  members (1) 
      -- CP-element group 415: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(415) is bound as output of CP function.
    -- CP-element group 416:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (1) 
      -- CP-element group 416: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(416) is bound as output of CP function.
    -- CP-element group 417:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	415 
    -- CP-element group 417: marked-predecessors 
    -- CP-element group 417: 	419 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	419 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/rr
      -- CP-element group 417: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/$entry
      -- 
    rr_1764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(417), ack => type_cast_842_inst_req_0); -- 
    concat_cp_element_group_417: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_417"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(415) & concat_CP_34_elements(419);
      gj_concat_cp_element_group_417 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(417), clk => clk, reset => reset); --
    end block;
    -- CP-element group 418:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: marked-predecessors 
    -- CP-element group 418: 	420 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	420 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/cr
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_start_
      -- 
    cr_1769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(418), ack => type_cast_842_inst_req_1); -- 
    concat_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(416) & concat_CP_34_elements(420);
      gj_concat_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419: marked-successors 
    -- CP-element group 419: 	417 
    -- CP-element group 419:  members (4) 
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_completed__ps
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/ra
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_completed_
      -- 
    ra_1765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_0, ack => concat_CP_34_elements(419)); -- 
    -- CP-element group 420:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	418 
    -- CP-element group 420: successors 
    -- CP-element group 420: marked-successors 
    -- CP-element group 420: 	418 
    -- CP-element group 420:  members (4) 
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_completed__ps
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/ca
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_completed_
      -- 
    ca_1770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_1, ack => concat_CP_34_elements(420)); -- 
    -- CP-element group 421:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: successors 
    -- CP-element group 421:  members (4) 
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_completed_
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_start_
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_completed__ps
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(421) is bound as output of CP function.
    -- CP-element group 422:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	424 
    -- CP-element group 422:  members (2) 
      -- CP-element group 422: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_start_
      -- CP-element group 422: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(422) is bound as output of CP function.
    -- CP-element group 423:  join  transition  bypass  pipeline-parent 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	424 
    -- CP-element group 423: successors 
    -- CP-element group 423:  members (1) 
      -- CP-element group 423: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_completed__ps
      -- 
    concat_CP_34_elements(423) <= concat_CP_34_elements(424);
    -- CP-element group 424:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	422 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	423 
    -- CP-element group 424:  members (1) 
      -- CP-element group 424: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_completed_
      -- 
    -- Element group concat_CP_34_elements(424) is a control-delay.
    cp_element_424_delay: control_delay_element  generic map(name => " 424_delay", delay_value => 1)  port map(req => concat_CP_34_elements(422), ack => concat_CP_34_elements(424), clk => clk, reset =>reset);
    -- CP-element group 425:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	388 
    -- CP-element group 425: marked-predecessors 
    -- CP-element group 425: 	427 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	427 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_sample_start_
      -- CP-element group 425: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/rr
      -- CP-element group 425: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/$entry
      -- 
    rr_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(425), ack => type_cast_847_inst_req_0); -- 
    concat_cp_element_group_425: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_425"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(388) & concat_CP_34_elements(427);
      gj_concat_cp_element_group_425 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(425), clk => clk, reset => reset); --
    end block;
    -- CP-element group 426:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	319 
    -- CP-element group 426: marked-predecessors 
    -- CP-element group 426: 	428 
    -- CP-element group 426: 	435 
    -- CP-element group 426: 	446 
    -- CP-element group 426: 	458 
    -- CP-element group 426: 	469 
    -- CP-element group 426: 	505 
    -- CP-element group 426: 	509 
    -- CP-element group 426: 	513 
    -- CP-element group 426: 	517 
    -- CP-element group 426: 	564 
    -- CP-element group 426: 	599 
    -- CP-element group 426: 	603 
    -- CP-element group 426: 	655 
    -- CP-element group 426: 	663 
    -- CP-element group 426: 	667 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	428 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/cr
      -- CP-element group 426: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/$entry
      -- CP-element group 426: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_update_start_
      -- 
    cr_1792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(426), ack => type_cast_847_inst_req_1); -- 
    concat_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(428) & concat_CP_34_elements(435) & concat_CP_34_elements(446) & concat_CP_34_elements(458) & concat_CP_34_elements(469) & concat_CP_34_elements(505) & concat_CP_34_elements(509) & concat_CP_34_elements(513) & concat_CP_34_elements(517) & concat_CP_34_elements(564) & concat_CP_34_elements(599) & concat_CP_34_elements(603) & concat_CP_34_elements(655) & concat_CP_34_elements(663) & concat_CP_34_elements(667);
      gj_concat_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	425 
    -- CP-element group 427: successors 
    -- CP-element group 427: marked-successors 
    -- CP-element group 427: 	384 
    -- CP-element group 427: 	425 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/ra
      -- CP-element group 427: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_sample_completed_
      -- CP-element group 427: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/$exit
      -- 
    ra_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_0, ack => concat_CP_34_elements(427)); -- 
    -- CP-element group 428:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	433 
    -- CP-element group 428: 	444 
    -- CP-element group 428: 	456 
    -- CP-element group 428: 	467 
    -- CP-element group 428: 	503 
    -- CP-element group 428: 	507 
    -- CP-element group 428: 	511 
    -- CP-element group 428: 	515 
    -- CP-element group 428: 	562 
    -- CP-element group 428: 	597 
    -- CP-element group 428: 	601 
    -- CP-element group 428: 	653 
    -- CP-element group 428: 	661 
    -- CP-element group 428: 	665 
    -- CP-element group 428: marked-successors 
    -- CP-element group 428: 	343 
    -- CP-element group 428: 	426 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_update_completed_
      -- CP-element group 428: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/$exit
      -- CP-element group 428: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/ca
      -- 
    ca_1793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_1, ack => concat_CP_34_elements(428)); -- 
    -- CP-element group 429:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	346 
    -- CP-element group 429: marked-predecessors 
    -- CP-element group 429: 	431 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	431 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/req
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_sample_start_
      -- 
    req_1801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(429), ack => W_add_inp1x_x1_866_delayed_1_0_864_inst_req_0); -- 
    concat_cp_element_group_429: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_429"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(346) & concat_CP_34_elements(431);
      gj_concat_cp_element_group_429 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(429), clk => clk, reset => reset); --
    end block;
    -- CP-element group 430:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: marked-predecessors 
    -- CP-element group 430: 	432 
    -- CP-element group 430: 	435 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	432 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/req
      -- CP-element group 430: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_update_start_
      -- CP-element group 430: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/$entry
      -- 
    req_1806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(430), ack => W_add_inp1x_x1_866_delayed_1_0_864_inst_req_1); -- 
    concat_cp_element_group_430: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_430"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(432) & concat_CP_34_elements(435);
      gj_concat_cp_element_group_430 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(430), clk => clk, reset => reset); --
    end block;
    -- CP-element group 431:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	429 
    -- CP-element group 431: successors 
    -- CP-element group 431: marked-successors 
    -- CP-element group 431: 	344 
    -- CP-element group 431: 	429 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/ack
      -- CP-element group 431: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_sample_completed_
      -- 
    ack_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_0, ack => concat_CP_34_elements(431)); -- 
    -- CP-element group 432:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	430 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432: marked-successors 
    -- CP-element group 432: 	430 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/ack
      -- CP-element group 432: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_update_completed_
      -- 
    ack_1807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_1, ack => concat_CP_34_elements(432)); -- 
    -- CP-element group 433:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	428 
    -- CP-element group 433: 	432 
    -- CP-element group 433: marked-predecessors 
    -- CP-element group 433: 	435 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	435 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_sample_start_
      -- CP-element group 433: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/$entry
      -- CP-element group 433: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/rr
      -- 
    rr_1815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(433), ack => type_cast_870_inst_req_0); -- 
    concat_cp_element_group_433: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_433"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(432) & concat_CP_34_elements(435);
      gj_concat_cp_element_group_433 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(433), clk => clk, reset => reset); --
    end block;
    -- CP-element group 434:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: marked-predecessors 
    -- CP-element group 434: 	436 
    -- CP-element group 434: 	440 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	436 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_update_start_
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/$entry
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/cr
      -- 
    cr_1820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(434), ack => type_cast_870_inst_req_1); -- 
    concat_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(436) & concat_CP_34_elements(440);
      gj_concat_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	433 
    -- CP-element group 435: successors 
    -- CP-element group 435: marked-successors 
    -- CP-element group 435: 	426 
    -- CP-element group 435: 	430 
    -- CP-element group 435: 	433 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_sample_completed_
      -- CP-element group 435: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/ra
      -- 
    ra_1816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_0, ack => concat_CP_34_elements(435)); -- 
    -- CP-element group 436:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	434 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	440 
    -- CP-element group 436: marked-successors 
    -- CP-element group 436: 	434 
    -- CP-element group 436:  members (16) 
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/$entry
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_update_completed_
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resized_1
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scaled_1
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_computed_1
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/ca
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/req
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/$entry
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/scale_rename_ack
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/scale_rename_req
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/$exit
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/$entry
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/index_resize_ack
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/index_resize_req
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/$exit
      -- 
    ca_1821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_1, ack => concat_CP_34_elements(436)); -- 
    req_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(436), ack => array_obj_ref_876_index_offset_req_0); -- 
    -- CP-element group 437:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	441 
    -- CP-element group 437: marked-predecessors 
    -- CP-element group 437: 	442 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	442 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/req
      -- CP-element group 437: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/$entry
      -- 
    req_1861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(437), ack => addr_of_877_final_reg_req_0); -- 
    concat_cp_element_group_437: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_437"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(441) & concat_CP_34_elements(442);
      gj_concat_cp_element_group_437 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(437), clk => clk, reset => reset); --
    end block;
    -- CP-element group 438:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	316 
    -- CP-element group 438: marked-predecessors 
    -- CP-element group 438: 	443 
    -- CP-element group 438: 	450 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	443 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/req
      -- CP-element group 438: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_update_start_
      -- CP-element group 438: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/$entry
      -- 
    req_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(438), ack => addr_of_877_final_reg_req_1); -- 
    concat_cp_element_group_438: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_438"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(443) & concat_CP_34_elements(450);
      gj_concat_cp_element_group_438 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(438), clk => clk, reset => reset); --
    end block;
    -- CP-element group 439:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	316 
    -- CP-element group 439: marked-predecessors 
    -- CP-element group 439: 	441 
    -- CP-element group 439: 	442 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	441 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/req
      -- CP-element group 439: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/$entry
      -- CP-element group 439: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_update_start
      -- 
    req_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(439), ack => array_obj_ref_876_index_offset_req_1); -- 
    concat_cp_element_group_439: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_439"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(441) & concat_CP_34_elements(442);
      gj_concat_cp_element_group_439 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(439), clk => clk, reset => reset); --
    end block;
    -- CP-element group 440:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	436 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	691 
    -- CP-element group 440: marked-successors 
    -- CP-element group 440: 	434 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/ack
      -- CP-element group 440: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/$exit
      -- CP-element group 440: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_sample_complete
      -- 
    ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_0, ack => concat_CP_34_elements(440)); -- 
    -- CP-element group 441:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	439 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	437 
    -- CP-element group 441: marked-successors 
    -- CP-element group 441: 	439 
    -- CP-element group 441:  members (8) 
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_offset_calculated
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_root_address_calculated
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/sum_rename_ack
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/sum_rename_req
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/$exit
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/$entry
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/ack
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/$exit
      -- 
    ack_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_1, ack => concat_CP_34_elements(441)); -- 
    -- CP-element group 442:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	437 
    -- CP-element group 442: successors 
    -- CP-element group 442: marked-successors 
    -- CP-element group 442: 	437 
    -- CP-element group 442: 	439 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_sample_completed_
      -- CP-element group 442: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/ack
      -- CP-element group 442: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/$exit
      -- 
    ack_1862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_0, ack => concat_CP_34_elements(442)); -- 
    -- CP-element group 443:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	438 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	448 
    -- CP-element group 443: marked-successors 
    -- CP-element group 443: 	438 
    -- CP-element group 443:  members (19) 
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_root_address_calculated
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/$entry
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/base_resize_ack
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/$entry
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_address_resized
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/root_register_req
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/sum_rename_req
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/sum_rename_ack
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/root_register_ack
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/$entry
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/base_resize_req
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_address_calculated
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_address_calculated
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/ack
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_update_completed_
      -- 
    ack_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_1, ack => concat_CP_34_elements(443)); -- 
    -- CP-element group 444:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	428 
    -- CP-element group 444: marked-predecessors 
    -- CP-element group 444: 	446 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	446 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/req
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/$entry
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_sample_start_
      -- 
    req_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(444), ack => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_0); -- 
    concat_cp_element_group_444: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_444"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(446);
      gj_concat_cp_element_group_444 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(444), clk => clk, reset => reset); --
    end block;
    -- CP-element group 445:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: marked-predecessors 
    -- CP-element group 445: 	447 
    -- CP-element group 445: 	450 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	447 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/req
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_update_start_
      -- 
    req_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_1); -- 
    concat_cp_element_group_445: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_445"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(447) & concat_CP_34_elements(450);
      gj_concat_cp_element_group_445 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(445), clk => clk, reset => reset); --
    end block;
    -- CP-element group 446:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	444 
    -- CP-element group 446: successors 
    -- CP-element group 446: marked-successors 
    -- CP-element group 446: 	426 
    -- CP-element group 446: 	444 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/ack
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/$exit
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_sample_completed_
      -- 
    ack_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_0, ack => concat_CP_34_elements(446)); -- 
    -- CP-element group 447:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	445 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447: marked-successors 
    -- CP-element group 447: 	445 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/ack
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/$exit
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_update_completed_
      -- 
    ack_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_1, ack => concat_CP_34_elements(447)); -- 
    -- CP-element group 448:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	443 
    -- CP-element group 448: 	447 
    -- CP-element group 448: marked-predecessors 
    -- CP-element group 448: 	450 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	450 
    -- CP-element group 448:  members (5) 
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/$entry
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/$entry
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/rr
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/$entry
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_sample_start_
      -- 
    rr_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(448), ack => ptr_deref_885_load_0_req_0); -- 
    concat_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(443) & concat_CP_34_elements(447) & concat_CP_34_elements(450);
      gj_concat_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: marked-predecessors 
    -- CP-element group 449: 	451 
    -- CP-element group 449: 	477 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	451 
    -- CP-element group 449:  members (5) 
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/$entry
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/cr
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_update_start_
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/$entry
      -- 
    cr_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(449), ack => ptr_deref_885_load_0_req_1); -- 
    concat_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(451) & concat_CP_34_elements(477);
      gj_concat_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	448 
    -- CP-element group 450: successors 
    -- CP-element group 450: marked-successors 
    -- CP-element group 450: 	438 
    -- CP-element group 450: 	445 
    -- CP-element group 450: 	448 
    -- CP-element group 450:  members (5) 
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/$exit
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/$exit
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/$exit
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/ra
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_sample_completed_
      -- 
    ra_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_885_load_0_ack_0, ack => concat_CP_34_elements(450)); -- 
    -- CP-element group 451:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	449 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	475 
    -- CP-element group 451: marked-successors 
    -- CP-element group 451: 	449 
    -- CP-element group 451:  members (9) 
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/$exit
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/ca
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/$exit
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/$exit
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/merge_req
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/merge_ack
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_update_completed_
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/$exit
      -- 
    ca_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_885_load_0_ack_1, ack => concat_CP_34_elements(451)); -- 
    -- CP-element group 452:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	327 
    -- CP-element group 452: marked-predecessors 
    -- CP-element group 452: 	454 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	454 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_sample_start_
      -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(452), ack => W_add_outx_x1_883_delayed_1_0_887_inst_req_0); -- 
    concat_cp_element_group_452: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_452"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(327) & concat_CP_34_elements(454);
      gj_concat_cp_element_group_452 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(452), clk => clk, reset => reset); --
    end block;
    -- CP-element group 453:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: marked-predecessors 
    -- CP-element group 453: 	455 
    -- CP-element group 453: 	458 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	455 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/$entry
      -- CP-element group 453: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/req
      -- CP-element group 453: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_update_start_
      -- 
    req_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(453), ack => W_add_outx_x1_883_delayed_1_0_887_inst_req_1); -- 
    concat_cp_element_group_453: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_453"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(455) & concat_CP_34_elements(458);
      gj_concat_cp_element_group_453 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(453), clk => clk, reset => reset); --
    end block;
    -- CP-element group 454:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	452 
    -- CP-element group 454: successors 
    -- CP-element group 454: marked-successors 
    -- CP-element group 454: 	452 
    -- CP-element group 454: 	323 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/ack
      -- CP-element group 454: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/$exit
      -- CP-element group 454: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_sample_completed_
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_883_delayed_1_0_887_inst_ack_0, ack => concat_CP_34_elements(454)); -- 
    -- CP-element group 455:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	453 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455: marked-successors 
    -- CP-element group 455: 	453 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/$exit
      -- CP-element group 455: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/ack
      -- CP-element group 455: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_update_completed_
      -- 
    ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_883_delayed_1_0_887_inst_ack_1, ack => concat_CP_34_elements(455)); -- 
    -- CP-element group 456:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	428 
    -- CP-element group 456: 	455 
    -- CP-element group 456: marked-predecessors 
    -- CP-element group 456: 	458 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	458 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_sample_start_
      -- CP-element group 456: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/rr
      -- CP-element group 456: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/$entry
      -- 
    rr_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(456), ack => type_cast_893_inst_req_0); -- 
    concat_cp_element_group_456: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_456"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(455) & concat_CP_34_elements(458);
      gj_concat_cp_element_group_456 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(456), clk => clk, reset => reset); --
    end block;
    -- CP-element group 457:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: marked-predecessors 
    -- CP-element group 457: 	459 
    -- CP-element group 457: 	463 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	459 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_update_start_
      -- CP-element group 457: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/cr
      -- CP-element group 457: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/$entry
      -- 
    cr_1958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(457), ack => type_cast_893_inst_req_1); -- 
    concat_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(459) & concat_CP_34_elements(463);
      gj_concat_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	456 
    -- CP-element group 458: successors 
    -- CP-element group 458: marked-successors 
    -- CP-element group 458: 	426 
    -- CP-element group 458: 	453 
    -- CP-element group 458: 	456 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/ra
      -- CP-element group 458: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/$exit
      -- 
    ra_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_893_inst_ack_0, ack => concat_CP_34_elements(458)); -- 
    -- CP-element group 459:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	457 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	463 
    -- CP-element group 459: marked-successors 
    -- CP-element group 459: 	457 
    -- CP-element group 459:  members (16) 
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/$entry
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/index_resize_req
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/index_resize_ack
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/$entry
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/req
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_computed_1
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scaled_1
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/ca
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resized_1
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/scale_rename_ack
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/scale_rename_req
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/$entry
      -- 
    ca_1959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_893_inst_ack_1, ack => concat_CP_34_elements(459)); -- 
    req_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(459), ack => array_obj_ref_899_index_offset_req_0); -- 
    -- CP-element group 460:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	464 
    -- CP-element group 460: marked-predecessors 
    -- CP-element group 460: 	465 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	465 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/$entry
      -- CP-element group 460: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/req
      -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(460), ack => addr_of_900_final_reg_req_0); -- 
    concat_cp_element_group_460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(464) & concat_CP_34_elements(465);
      gj_concat_cp_element_group_460 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(460), clk => clk, reset => reset); --
    end block;
    -- CP-element group 461:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	316 
    -- CP-element group 461: marked-predecessors 
    -- CP-element group 461: 	466 
    -- CP-element group 461: 	473 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	466 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_update_start_
      -- CP-element group 461: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/req
      -- CP-element group 461: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/$entry
      -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(461), ack => addr_of_900_final_reg_req_1); -- 
    concat_cp_element_group_461: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_461"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(466) & concat_CP_34_elements(473);
      gj_concat_cp_element_group_461 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(461), clk => clk, reset => reset); --
    end block;
    -- CP-element group 462:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	316 
    -- CP-element group 462: marked-predecessors 
    -- CP-element group 462: 	464 
    -- CP-element group 462: 	465 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	464 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_update_start
      -- CP-element group 462: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/req
      -- CP-element group 462: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/$entry
      -- 
    req_1989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(462), ack => array_obj_ref_899_index_offset_req_1); -- 
    concat_cp_element_group_462: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_462"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(464) & concat_CP_34_elements(465);
      gj_concat_cp_element_group_462 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(462), clk => clk, reset => reset); --
    end block;
    -- CP-element group 463:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	459 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	691 
    -- CP-element group 463: marked-successors 
    -- CP-element group 463: 	457 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_sample_complete
      -- CP-element group 463: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/$exit
      -- CP-element group 463: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/ack
      -- 
    ack_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_899_index_offset_ack_0, ack => concat_CP_34_elements(463)); -- 
    -- CP-element group 464:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	460 
    -- CP-element group 464: marked-successors 
    -- CP-element group 464: 	462 
    -- CP-element group 464:  members (8) 
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/sum_rename_req
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/sum_rename_ack
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/$entry
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/$exit
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_offset_calculated
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_root_address_calculated
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/ack
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/$exit
      -- 
    ack_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_899_index_offset_ack_1, ack => concat_CP_34_elements(464)); -- 
    -- CP-element group 465:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	460 
    -- CP-element group 465: successors 
    -- CP-element group 465: marked-successors 
    -- CP-element group 465: 	460 
    -- CP-element group 465: 	462 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_sample_completed_
      -- CP-element group 465: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/ack
      -- CP-element group 465: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/$exit
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_900_final_reg_ack_0, ack => concat_CP_34_elements(465)); -- 
    -- CP-element group 466:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	461 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	471 
    -- CP-element group 466: marked-successors 
    -- CP-element group 466: 	461 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_update_completed_
      -- CP-element group 466: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/ack
      -- CP-element group 466: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/$exit
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_900_final_reg_ack_1, ack => concat_CP_34_elements(466)); -- 
    -- CP-element group 467:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	428 
    -- CP-element group 467: marked-predecessors 
    -- CP-element group 467: 	469 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	469 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_sample_start_
      -- CP-element group 467: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/req
      -- CP-element group 467: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/$entry
      -- 
    req_2013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(467), ack => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_0); -- 
    concat_cp_element_group_467: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_467"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(469);
      gj_concat_cp_element_group_467 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(467), clk => clk, reset => reset); --
    end block;
    -- CP-element group 468:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: marked-predecessors 
    -- CP-element group 468: 	470 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	470 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_update_start_
      -- CP-element group 468: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/req
      -- CP-element group 468: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/$entry
      -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(468), ack => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_1); -- 
    concat_cp_element_group_468: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_468"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(470);
      gj_concat_cp_element_group_468 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(468), clk => clk, reset => reset); --
    end block;
    -- CP-element group 469:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	467 
    -- CP-element group 469: successors 
    -- CP-element group 469: marked-successors 
    -- CP-element group 469: 	426 
    -- CP-element group 469: 	467 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_sample_completed_
      -- CP-element group 469: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/ack
      -- CP-element group 469: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/$exit
      -- 
    ack_2014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_0, ack => concat_CP_34_elements(469)); -- 
    -- CP-element group 470:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	468 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	691 
    -- CP-element group 470: marked-successors 
    -- CP-element group 470: 	468 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_update_completed_
      -- CP-element group 470: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/ack
      -- CP-element group 470: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/$exit
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_1, ack => concat_CP_34_elements(470)); -- 
    -- CP-element group 471:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	466 
    -- CP-element group 471: marked-predecessors 
    -- CP-element group 471: 	473 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	473 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_sample_start_
      -- CP-element group 471: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/req
      -- CP-element group 471: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/$entry
      -- 
    req_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(471), ack => W_arrayidx245_894_delayed_6_0_905_inst_req_0); -- 
    concat_cp_element_group_471: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_471"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(466) & concat_CP_34_elements(473);
      gj_concat_cp_element_group_471 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(471), clk => clk, reset => reset); --
    end block;
    -- CP-element group 472:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: marked-predecessors 
    -- CP-element group 472: 	474 
    -- CP-element group 472: 	477 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	474 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/req
      -- CP-element group 472: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/$entry
      -- CP-element group 472: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_update_start_
      -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(472), ack => W_arrayidx245_894_delayed_6_0_905_inst_req_1); -- 
    concat_cp_element_group_472: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_472"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(474) & concat_CP_34_elements(477);
      gj_concat_cp_element_group_472 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(472), clk => clk, reset => reset); --
    end block;
    -- CP-element group 473:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	471 
    -- CP-element group 473: successors 
    -- CP-element group 473: marked-successors 
    -- CP-element group 473: 	461 
    -- CP-element group 473: 	471 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_sample_completed_
      -- CP-element group 473: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/ack
      -- CP-element group 473: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/$exit
      -- 
    ack_2028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx245_894_delayed_6_0_905_inst_ack_0, ack => concat_CP_34_elements(473)); -- 
    -- CP-element group 474:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	472 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474: marked-successors 
    -- CP-element group 474: 	472 
    -- CP-element group 474:  members (19) 
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/root_register_req
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_address_resized
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/$entry
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/$exit
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/base_resize_req
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_root_address_calculated
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/$exit
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/$entry
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/$entry
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/$exit
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_address_calculated
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/sum_rename_ack
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_address_calculated
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/ack
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/$exit
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/sum_rename_req
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/base_resize_ack
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/root_register_ack
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_update_completed_
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx245_894_delayed_6_0_905_inst_ack_1, ack => concat_CP_34_elements(474)); -- 
    -- CP-element group 475:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	451 
    -- CP-element group 475: 	474 
    -- CP-element group 475: marked-predecessors 
    -- CP-element group 475: 	477 
    -- CP-element group 475: 	587 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	477 
    -- CP-element group 475:  members (9) 
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/split_req
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/$entry
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/$exit
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/$entry
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/$entry
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/rr
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/split_ack
      -- 
    rr_2071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(475), ack => ptr_deref_910_store_0_req_0); -- 
    concat_cp_element_group_475: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_475"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(451) & concat_CP_34_elements(474) & concat_CP_34_elements(477) & concat_CP_34_elements(587);
      gj_concat_cp_element_group_475 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(475), clk => clk, reset => reset); --
    end block;
    -- CP-element group 476:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: marked-predecessors 
    -- CP-element group 476: 	478 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	478 
    -- CP-element group 476:  members (5) 
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_update_start_
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/cr
      -- 
    cr_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(476), ack => ptr_deref_910_store_0_req_1); -- 
    concat_cp_element_group_476: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_476"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(478);
      gj_concat_cp_element_group_476 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(476), clk => clk, reset => reset); --
    end block;
    -- CP-element group 477:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	475 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	690 
    -- CP-element group 477: marked-successors 
    -- CP-element group 477: 	449 
    -- CP-element group 477: 	472 
    -- CP-element group 477: 	475 
    -- CP-element group 477:  members (5) 
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_sample_completed_
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/$exit
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/$exit
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/$exit
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/ra
      -- 
    ra_2072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_910_store_0_ack_0, ack => concat_CP_34_elements(477)); -- 
    -- CP-element group 478:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	476 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	691 
    -- CP-element group 478: marked-successors 
    -- CP-element group 478: 	476 
    -- CP-element group 478:  members (5) 
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_update_completed_
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/$exit
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/$exit
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/$exit
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/ca
      -- 
    ca_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_910_store_0_ack_1, ack => concat_CP_34_elements(478)); -- 
    -- CP-element group 479:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	388 
    -- CP-element group 479: marked-predecessors 
    -- CP-element group 479: 	481 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	481 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_sample_start_
      -- CP-element group 479: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/$entry
      -- CP-element group 479: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/req
      -- 
    req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(479), ack => W_count_inp1x_x1_900_delayed_1_0_913_inst_req_0); -- 
    concat_cp_element_group_479: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_479"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(388) & concat_CP_34_elements(481);
      gj_concat_cp_element_group_479 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(479), clk => clk, reset => reset); --
    end block;
    -- CP-element group 480:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: marked-predecessors 
    -- CP-element group 480: 	482 
    -- CP-element group 480: 	505 
    -- CP-element group 480: 	663 
    -- CP-element group 480: 	667 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	482 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_update_start_
      -- CP-element group 480: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/$entry
      -- CP-element group 480: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/req
      -- 
    req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(480), ack => W_count_inp1x_x1_900_delayed_1_0_913_inst_req_1); -- 
    concat_cp_element_group_480: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_480"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(482) & concat_CP_34_elements(505) & concat_CP_34_elements(663) & concat_CP_34_elements(667);
      gj_concat_cp_element_group_480 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(480), clk => clk, reset => reset); --
    end block;
    -- CP-element group 481:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	479 
    -- CP-element group 481: successors 
    -- CP-element group 481: marked-successors 
    -- CP-element group 481: 	384 
    -- CP-element group 481: 	479 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_sample_completed_
      -- CP-element group 481: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/$exit
      -- CP-element group 481: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/ack
      -- 
    ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_0, ack => concat_CP_34_elements(481)); -- 
    -- CP-element group 482:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	480 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	503 
    -- CP-element group 482: 	661 
    -- CP-element group 482: 	665 
    -- CP-element group 482: marked-successors 
    -- CP-element group 482: 	480 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_update_completed_
      -- CP-element group 482: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/$exit
      -- CP-element group 482: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/ack
      -- 
    ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_1, ack => concat_CP_34_elements(482)); -- 
    -- CP-element group 483:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	346 
    -- CP-element group 483: marked-predecessors 
    -- CP-element group 483: 	485 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	485 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/req
      -- 
    req_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(483), ack => W_add_inp1x_x1_907_delayed_1_0_923_inst_req_0); -- 
    concat_cp_element_group_483: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_483"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(346) & concat_CP_34_elements(485);
      gj_concat_cp_element_group_483 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(483), clk => clk, reset => reset); --
    end block;
    -- CP-element group 484:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	319 
    -- CP-element group 484: marked-predecessors 
    -- CP-element group 484: 	486 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	486 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_update_start_
      -- CP-element group 484: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/req
      -- 
    req_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(484), ack => W_add_inp1x_x1_907_delayed_1_0_923_inst_req_1); -- 
    concat_cp_element_group_484: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_484"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(486);
      gj_concat_cp_element_group_484 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(484), clk => clk, reset => reset); --
    end block;
    -- CP-element group 485:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	483 
    -- CP-element group 485: successors 
    -- CP-element group 485: marked-successors 
    -- CP-element group 485: 	344 
    -- CP-element group 485: 	483 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_sample_completed_
      -- CP-element group 485: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/ack
      -- 
    ack_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_0, ack => concat_CP_34_elements(485)); -- 
    -- CP-element group 486:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	484 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	691 
    -- CP-element group 486: marked-successors 
    -- CP-element group 486: 	343 
    -- CP-element group 486: 	484 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_update_completed_
      -- CP-element group 486: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/ack
      -- 
    ack_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_1, ack => concat_CP_34_elements(486)); -- 
    -- CP-element group 487:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	327 
    -- CP-element group 487: marked-predecessors 
    -- CP-element group 487: 	489 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	489 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_sample_start_
      -- CP-element group 487: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/$entry
      -- CP-element group 487: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/req
      -- 
    req_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(487), ack => W_add_outx_x1_914_delayed_1_0_933_inst_req_0); -- 
    concat_cp_element_group_487: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_487"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(327) & concat_CP_34_elements(489);
      gj_concat_cp_element_group_487 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(487), clk => clk, reset => reset); --
    end block;
    -- CP-element group 488:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: marked-predecessors 
    -- CP-element group 488: 	490 
    -- CP-element group 488: 	564 
    -- CP-element group 488: 	599 
    -- CP-element group 488: 	603 
    -- CP-element group 488: 	655 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	490 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_update_start_
      -- CP-element group 488: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/req
      -- 
    req_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(488), ack => W_add_outx_x1_914_delayed_1_0_933_inst_req_1); -- 
    concat_cp_element_group_488: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_488"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(490) & concat_CP_34_elements(564) & concat_CP_34_elements(599) & concat_CP_34_elements(603) & concat_CP_34_elements(655);
      gj_concat_cp_element_group_488 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(488), clk => clk, reset => reset); --
    end block;
    -- CP-element group 489:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	487 
    -- CP-element group 489: successors 
    -- CP-element group 489: marked-successors 
    -- CP-element group 489: 	487 
    -- CP-element group 489: 	323 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_sample_completed_
      -- CP-element group 489: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/$exit
      -- CP-element group 489: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/ack
      -- 
    ack_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_914_delayed_1_0_933_inst_ack_0, ack => concat_CP_34_elements(489)); -- 
    -- CP-element group 490:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	488 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	562 
    -- CP-element group 490: 	597 
    -- CP-element group 490: 	601 
    -- CP-element group 490: 	653 
    -- CP-element group 490: marked-successors 
    -- CP-element group 490: 	488 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_update_completed_
      -- CP-element group 490: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/$exit
      -- CP-element group 490: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/ack
      -- 
    ack_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_914_delayed_1_0_933_inst_ack_1, ack => concat_CP_34_elements(490)); -- 
    -- CP-element group 491:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	327 
    -- CP-element group 491: marked-predecessors 
    -- CP-element group 491: 	493 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	493 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_sample_start_
      -- CP-element group 491: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/$entry
      -- CP-element group 491: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/rr
      -- 
    rr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(491), ack => type_cast_953_inst_req_0); -- 
    concat_cp_element_group_491: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_491"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(327) & concat_CP_34_elements(493);
      gj_concat_cp_element_group_491 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(491), clk => clk, reset => reset); --
    end block;
    -- CP-element group 492:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: marked-predecessors 
    -- CP-element group 492: 	494 
    -- CP-element group 492: 	564 
    -- CP-element group 492: 	599 
    -- CP-element group 492: 	603 
    -- CP-element group 492: 	655 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	494 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_update_start_
      -- CP-element group 492: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/$entry
      -- CP-element group 492: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/cr
      -- 
    cr_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(492), ack => type_cast_953_inst_req_1); -- 
    concat_cp_element_group_492: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_492"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(494) & concat_CP_34_elements(564) & concat_CP_34_elements(599) & concat_CP_34_elements(603) & concat_CP_34_elements(655);
      gj_concat_cp_element_group_492 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(492), clk => clk, reset => reset); --
    end block;
    -- CP-element group 493:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	491 
    -- CP-element group 493: successors 
    -- CP-element group 493: marked-successors 
    -- CP-element group 493: 	491 
    -- CP-element group 493: 	323 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_sample_completed_
      -- CP-element group 493: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/$exit
      -- CP-element group 493: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/ra
      -- 
    ra_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_953_inst_ack_0, ack => concat_CP_34_elements(493)); -- 
    -- CP-element group 494:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	492 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	562 
    -- CP-element group 494: 	597 
    -- CP-element group 494: 	601 
    -- CP-element group 494: 	653 
    -- CP-element group 494: marked-successors 
    -- CP-element group 494: 	492 
    -- CP-element group 494:  members (3) 
      -- CP-element group 494: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_update_completed_
      -- CP-element group 494: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/$exit
      -- CP-element group 494: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/ca
      -- 
    ca_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_953_inst_ack_1, ack => concat_CP_34_elements(494)); -- 
    -- CP-element group 495:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	346 
    -- CP-element group 495: marked-predecessors 
    -- CP-element group 495: 	497 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	497 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_sample_start_
      -- CP-element group 495: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/$entry
      -- CP-element group 495: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/rr
      -- 
    rr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(495), ack => type_cast_968_inst_req_0); -- 
    concat_cp_element_group_495: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_495"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(346) & concat_CP_34_elements(497);
      gj_concat_cp_element_group_495 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(495), clk => clk, reset => reset); --
    end block;
    -- CP-element group 496:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	319 
    -- CP-element group 496: marked-predecessors 
    -- CP-element group 496: 	498 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	498 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_update_start_
      -- CP-element group 496: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/cr
      -- 
    cr_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(496), ack => type_cast_968_inst_req_1); -- 
    concat_cp_element_group_496: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_496"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(498);
      gj_concat_cp_element_group_496 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 497:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	495 
    -- CP-element group 497: successors 
    -- CP-element group 497: marked-successors 
    -- CP-element group 497: 	344 
    -- CP-element group 497: 	495 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_sample_completed_
      -- CP-element group 497: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/$exit
      -- CP-element group 497: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/ra
      -- 
    ra_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_0, ack => concat_CP_34_elements(497)); -- 
    -- CP-element group 498:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	496 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	691 
    -- CP-element group 498: marked-successors 
    -- CP-element group 498: 	343 
    -- CP-element group 498: 	496 
    -- CP-element group 498:  members (3) 
      -- CP-element group 498: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_update_completed_
      -- CP-element group 498: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/$exit
      -- CP-element group 498: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/ca
      -- 
    ca_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_1, ack => concat_CP_34_elements(498)); -- 
    -- CP-element group 499:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	388 
    -- CP-element group 499: marked-predecessors 
    -- CP-element group 499: 	501 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	501 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_sample_start_
      -- CP-element group 499: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/rr
      -- 
    rr_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(499), ack => type_cast_983_inst_req_0); -- 
    concat_cp_element_group_499: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_499"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(388) & concat_CP_34_elements(501);
      gj_concat_cp_element_group_499 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(499), clk => clk, reset => reset); --
    end block;
    -- CP-element group 500:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: marked-predecessors 
    -- CP-element group 500: 	502 
    -- CP-element group 500: 	505 
    -- CP-element group 500: 	663 
    -- CP-element group 500: 	667 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	502 
    -- CP-element group 500:  members (3) 
      -- CP-element group 500: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_update_start_
      -- CP-element group 500: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/$entry
      -- CP-element group 500: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/cr
      -- 
    cr_2166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(500), ack => type_cast_983_inst_req_1); -- 
    concat_cp_element_group_500: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_500"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(502) & concat_CP_34_elements(505) & concat_CP_34_elements(663) & concat_CP_34_elements(667);
      gj_concat_cp_element_group_500 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(500), clk => clk, reset => reset); --
    end block;
    -- CP-element group 501:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	499 
    -- CP-element group 501: successors 
    -- CP-element group 501: marked-successors 
    -- CP-element group 501: 	384 
    -- CP-element group 501: 	499 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_sample_completed_
      -- CP-element group 501: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/$exit
      -- CP-element group 501: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/ra
      -- 
    ra_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_983_inst_ack_0, ack => concat_CP_34_elements(501)); -- 
    -- CP-element group 502:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	500 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	503 
    -- CP-element group 502: 	661 
    -- CP-element group 502: 	665 
    -- CP-element group 502: marked-successors 
    -- CP-element group 502: 	500 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_update_completed_
      -- CP-element group 502: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/$exit
      -- CP-element group 502: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/ca
      -- 
    ca_2167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_983_inst_ack_1, ack => concat_CP_34_elements(502)); -- 
    -- CP-element group 503:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	428 
    -- CP-element group 503: 	482 
    -- CP-element group 503: 	502 
    -- CP-element group 503: marked-predecessors 
    -- CP-element group 503: 	505 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	505 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_sample_start_
      -- CP-element group 503: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/rr
      -- 
    rr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(503), ack => type_cast_999_inst_req_0); -- 
    concat_cp_element_group_503: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_503"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(482) & concat_CP_34_elements(502) & concat_CP_34_elements(505);
      gj_concat_cp_element_group_503 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(503), clk => clk, reset => reset); --
    end block;
    -- CP-element group 504:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: marked-predecessors 
    -- CP-element group 504: 	506 
    -- CP-element group 504: 	525 
    -- CP-element group 504: 	529 
    -- CP-element group 504: 	533 
    -- CP-element group 504: 	537 
    -- CP-element group 504: 	643 
    -- CP-element group 504: 	659 
    -- CP-element group 504: 	671 
    -- CP-element group 504: 	683 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	506 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_update_start_
      -- CP-element group 504: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/cr
      -- 
    cr_2180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(504), ack => type_cast_999_inst_req_1); -- 
    concat_cp_element_group_504: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_504"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(525) & concat_CP_34_elements(529) & concat_CP_34_elements(533) & concat_CP_34_elements(537) & concat_CP_34_elements(643) & concat_CP_34_elements(659) & concat_CP_34_elements(671) & concat_CP_34_elements(683);
      gj_concat_cp_element_group_504 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(504), clk => clk, reset => reset); --
    end block;
    -- CP-element group 505:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	503 
    -- CP-element group 505: successors 
    -- CP-element group 505: marked-successors 
    -- CP-element group 505: 	426 
    -- CP-element group 505: 	480 
    -- CP-element group 505: 	500 
    -- CP-element group 505: 	503 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_sample_completed_
      -- CP-element group 505: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/$exit
      -- CP-element group 505: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/ra
      -- 
    ra_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_999_inst_ack_0, ack => concat_CP_34_elements(505)); -- 
    -- CP-element group 506:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	504 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	523 
    -- CP-element group 506: 	527 
    -- CP-element group 506: 	531 
    -- CP-element group 506: 	535 
    -- CP-element group 506: 	641 
    -- CP-element group 506: 	657 
    -- CP-element group 506: 	669 
    -- CP-element group 506: 	681 
    -- CP-element group 506: marked-successors 
    -- CP-element group 506: 	504 
    -- CP-element group 506:  members (3) 
      -- CP-element group 506: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_update_completed_
      -- CP-element group 506: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/$exit
      -- CP-element group 506: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/ca
      -- 
    ca_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_999_inst_ack_1, ack => concat_CP_34_elements(506)); -- 
    -- CP-element group 507:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	428 
    -- CP-element group 507: marked-predecessors 
    -- CP-element group 507: 	509 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	509 
    -- CP-element group 507:  members (3) 
      -- CP-element group 507: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/req
      -- 
    req_2189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(507), ack => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_0); -- 
    concat_cp_element_group_507: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_507"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(509);
      gj_concat_cp_element_group_507 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(507), clk => clk, reset => reset); --
    end block;
    -- CP-element group 508:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: marked-predecessors 
    -- CP-element group 508: 	510 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	510 
    -- CP-element group 508:  members (3) 
      -- CP-element group 508: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_update_start_
      -- CP-element group 508: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/$entry
      -- CP-element group 508: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/req
      -- 
    req_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(508), ack => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_1); -- 
    concat_cp_element_group_508: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_508"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(510);
      gj_concat_cp_element_group_508 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(508), clk => clk, reset => reset); --
    end block;
    -- CP-element group 509:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	507 
    -- CP-element group 509: successors 
    -- CP-element group 509: marked-successors 
    -- CP-element group 509: 	426 
    -- CP-element group 509: 	507 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_sample_completed_
      -- CP-element group 509: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/$exit
      -- CP-element group 509: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/ack
      -- 
    ack_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_0, ack => concat_CP_34_elements(509)); -- 
    -- CP-element group 510:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	508 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	691 
    -- CP-element group 510: marked-successors 
    -- CP-element group 510: 	508 
    -- CP-element group 510:  members (3) 
      -- CP-element group 510: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_update_completed_
      -- CP-element group 510: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/$exit
      -- CP-element group 510: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/ack
      -- 
    ack_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_1, ack => concat_CP_34_elements(510)); -- 
    -- CP-element group 511:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	428 
    -- CP-element group 511: marked-predecessors 
    -- CP-element group 511: 	513 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	513 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_sample_start_
      -- CP-element group 511: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/$entry
      -- CP-element group 511: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/req
      -- 
    req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(511), ack => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_0); -- 
    concat_cp_element_group_511: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_511"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(513);
      gj_concat_cp_element_group_511 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(511), clk => clk, reset => reset); --
    end block;
    -- CP-element group 512:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: marked-predecessors 
    -- CP-element group 512: 	514 
    -- CP-element group 512: 	525 
    -- CP-element group 512: 	529 
    -- CP-element group 512: 	533 
    -- CP-element group 512: 	537 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	514 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_update_start_
      -- CP-element group 512: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/$entry
      -- CP-element group 512: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/req
      -- 
    req_2208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(512), ack => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_1); -- 
    concat_cp_element_group_512: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_512"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(514) & concat_CP_34_elements(525) & concat_CP_34_elements(529) & concat_CP_34_elements(533) & concat_CP_34_elements(537);
      gj_concat_cp_element_group_512 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(512), clk => clk, reset => reset); --
    end block;
    -- CP-element group 513:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	511 
    -- CP-element group 513: successors 
    -- CP-element group 513: marked-successors 
    -- CP-element group 513: 	426 
    -- CP-element group 513: 	511 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_sample_completed_
      -- CP-element group 513: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/$exit
      -- CP-element group 513: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/ack
      -- 
    ack_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_0, ack => concat_CP_34_elements(513)); -- 
    -- CP-element group 514:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	512 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	523 
    -- CP-element group 514: 	527 
    -- CP-element group 514: 	531 
    -- CP-element group 514: 	535 
    -- CP-element group 514: marked-successors 
    -- CP-element group 514: 	512 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_update_completed_
      -- CP-element group 514: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/$exit
      -- CP-element group 514: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/ack
      -- 
    ack_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_1, ack => concat_CP_34_elements(514)); -- 
    -- CP-element group 515:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	428 
    -- CP-element group 515: marked-predecessors 
    -- CP-element group 515: 	517 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	517 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_sample_start_
      -- CP-element group 515: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/$entry
      -- CP-element group 515: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/req
      -- 
    req_2217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(515), ack => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_0); -- 
    concat_cp_element_group_515: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_515"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(517);
      gj_concat_cp_element_group_515 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(515), clk => clk, reset => reset); --
    end block;
    -- CP-element group 516:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: marked-predecessors 
    -- CP-element group 516: 	518 
    -- CP-element group 516: 	643 
    -- CP-element group 516: 	659 
    -- CP-element group 516: 	671 
    -- CP-element group 516: 	683 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	518 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_update_start_
      -- CP-element group 516: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/$entry
      -- CP-element group 516: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/req
      -- 
    req_2222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(516), ack => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_1); -- 
    concat_cp_element_group_516: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_516"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(518) & concat_CP_34_elements(643) & concat_CP_34_elements(659) & concat_CP_34_elements(671) & concat_CP_34_elements(683);
      gj_concat_cp_element_group_516 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(516), clk => clk, reset => reset); --
    end block;
    -- CP-element group 517:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	515 
    -- CP-element group 517: successors 
    -- CP-element group 517: marked-successors 
    -- CP-element group 517: 	426 
    -- CP-element group 517: 	515 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_sample_completed_
      -- CP-element group 517: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/$exit
      -- CP-element group 517: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/ack
      -- 
    ack_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_0, ack => concat_CP_34_elements(517)); -- 
    -- CP-element group 518:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	516 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	641 
    -- CP-element group 518: 	657 
    -- CP-element group 518: 	669 
    -- CP-element group 518: 	681 
    -- CP-element group 518: marked-successors 
    -- CP-element group 518: 	516 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_update_completed_
      -- CP-element group 518: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/$exit
      -- CP-element group 518: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/ack
      -- 
    ack_2223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_1, ack => concat_CP_34_elements(518)); -- 
    -- CP-element group 519:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	409 
    -- CP-element group 519: marked-predecessors 
    -- CP-element group 519: 	521 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	521 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_sample_start_
      -- CP-element group 519: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/$entry
      -- CP-element group 519: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/req
      -- 
    req_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(519), ack => W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_0); -- 
    concat_cp_element_group_519: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_519"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(409) & concat_CP_34_elements(521);
      gj_concat_cp_element_group_519 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(519), clk => clk, reset => reset); --
    end block;
    -- CP-element group 520:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: marked-predecessors 
    -- CP-element group 520: 	522 
    -- CP-element group 520: 	525 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	522 
    -- CP-element group 520:  members (3) 
      -- CP-element group 520: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_update_start_
      -- CP-element group 520: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/req
      -- 
    req_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(520), ack => W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_1); -- 
    concat_cp_element_group_520: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_520"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(522) & concat_CP_34_elements(525);
      gj_concat_cp_element_group_520 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(520), clk => clk, reset => reset); --
    end block;
    -- CP-element group 521:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	519 
    -- CP-element group 521: successors 
    -- CP-element group 521: marked-successors 
    -- CP-element group 521: 	405 
    -- CP-element group 521: 	519 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_sample_completed_
      -- CP-element group 521: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/$exit
      -- CP-element group 521: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/ack
      -- 
    ack_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_0, ack => concat_CP_34_elements(521)); -- 
    -- CP-element group 522:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	520 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	523 
    -- CP-element group 522: marked-successors 
    -- CP-element group 522: 	520 
    -- CP-element group 522:  members (3) 
      -- CP-element group 522: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_update_completed_
      -- CP-element group 522: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/$exit
      -- CP-element group 522: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/ack
      -- 
    ack_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 522_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_1, ack => concat_CP_34_elements(522)); -- 
    -- CP-element group 523:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	506 
    -- CP-element group 523: 	514 
    -- CP-element group 523: 	522 
    -- CP-element group 523: marked-predecessors 
    -- CP-element group 523: 	525 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	525 
    -- CP-element group 523:  members (3) 
      -- CP-element group 523: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_sample_start_
      -- CP-element group 523: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/$entry
      -- CP-element group 523: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/rr
      -- 
    rr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(523), ack => type_cast_1036_inst_req_0); -- 
    concat_cp_element_group_523: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_523"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(514) & concat_CP_34_elements(522) & concat_CP_34_elements(525);
      gj_concat_cp_element_group_523 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(523), clk => clk, reset => reset); --
    end block;
    -- CP-element group 524:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: marked-predecessors 
    -- CP-element group 524: 	526 
    -- CP-element group 524: 	545 
    -- CP-element group 524: 	556 
    -- CP-element group 524: 	568 
    -- CP-element group 524: 	579 
    -- CP-element group 524: 	615 
    -- CP-element group 524: 	619 
    -- CP-element group 524: 	623 
    -- CP-element group 524: 	627 
    -- CP-element group 524: 	631 
    -- CP-element group 524: 	635 
    -- CP-element group 524: 	647 
    -- CP-element group 524: 	651 
    -- CP-element group 524: 	675 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	526 
    -- CP-element group 524:  members (3) 
      -- CP-element group 524: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_update_start_
      -- CP-element group 524: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/$entry
      -- CP-element group 524: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/cr
      -- 
    cr_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(524), ack => type_cast_1036_inst_req_1); -- 
    concat_cp_element_group_524: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_524"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(545) & concat_CP_34_elements(556) & concat_CP_34_elements(568) & concat_CP_34_elements(579) & concat_CP_34_elements(615) & concat_CP_34_elements(619) & concat_CP_34_elements(623) & concat_CP_34_elements(627) & concat_CP_34_elements(631) & concat_CP_34_elements(635) & concat_CP_34_elements(647) & concat_CP_34_elements(651) & concat_CP_34_elements(675);
      gj_concat_cp_element_group_524 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(524), clk => clk, reset => reset); --
    end block;
    -- CP-element group 525:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	523 
    -- CP-element group 525: successors 
    -- CP-element group 525: marked-successors 
    -- CP-element group 525: 	504 
    -- CP-element group 525: 	512 
    -- CP-element group 525: 	520 
    -- CP-element group 525: 	523 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_sample_completed_
      -- CP-element group 525: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/$exit
      -- CP-element group 525: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/ra
      -- 
    ra_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1036_inst_ack_0, ack => concat_CP_34_elements(525)); -- 
    -- CP-element group 526:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	524 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	543 
    -- CP-element group 526: 	554 
    -- CP-element group 526: 	566 
    -- CP-element group 526: 	577 
    -- CP-element group 526: 	613 
    -- CP-element group 526: 	617 
    -- CP-element group 526: 	621 
    -- CP-element group 526: 	625 
    -- CP-element group 526: 	629 
    -- CP-element group 526: 	633 
    -- CP-element group 526: 	645 
    -- CP-element group 526: 	649 
    -- CP-element group 526: 	673 
    -- CP-element group 526: marked-successors 
    -- CP-element group 526: 	524 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_update_completed_
      -- CP-element group 526: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/$exit
      -- CP-element group 526: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/ca
      -- 
    ca_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 526_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1036_inst_ack_1, ack => concat_CP_34_elements(526)); -- 
    -- CP-element group 527:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	506 
    -- CP-element group 527: 	514 
    -- CP-element group 527: marked-predecessors 
    -- CP-element group 527: 	529 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	529 
    -- CP-element group 527:  members (3) 
      -- CP-element group 527: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_sample_start_
      -- CP-element group 527: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/$entry
      -- CP-element group 527: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/req
      -- 
    req_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(527), ack => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_0); -- 
    concat_cp_element_group_527: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_527"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(514) & concat_CP_34_elements(529);
      gj_concat_cp_element_group_527 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(527), clk => clk, reset => reset); --
    end block;
    -- CP-element group 528:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: marked-predecessors 
    -- CP-element group 528: 	530 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	530 
    -- CP-element group 528:  members (3) 
      -- CP-element group 528: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_update_start_
      -- CP-element group 528: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/req
      -- 
    req_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(528), ack => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_1); -- 
    concat_cp_element_group_528: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_528"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(530);
      gj_concat_cp_element_group_528 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(528), clk => clk, reset => reset); --
    end block;
    -- CP-element group 529:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	527 
    -- CP-element group 529: successors 
    -- CP-element group 529: marked-successors 
    -- CP-element group 529: 	504 
    -- CP-element group 529: 	512 
    -- CP-element group 529: 	527 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_sample_completed_
      -- CP-element group 529: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/$exit
      -- CP-element group 529: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/ack
      -- 
    ack_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 529_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_0, ack => concat_CP_34_elements(529)); -- 
    -- CP-element group 530:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	528 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	691 
    -- CP-element group 530: marked-successors 
    -- CP-element group 530: 	528 
    -- CP-element group 530:  members (3) 
      -- CP-element group 530: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_update_completed_
      -- CP-element group 530: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/$exit
      -- CP-element group 530: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/ack
      -- 
    ack_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_1, ack => concat_CP_34_elements(530)); -- 
    -- CP-element group 531:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	506 
    -- CP-element group 531: 	514 
    -- CP-element group 531: marked-predecessors 
    -- CP-element group 531: 	533 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	533 
    -- CP-element group 531:  members (3) 
      -- CP-element group 531: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_sample_start_
      -- CP-element group 531: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/$entry
      -- CP-element group 531: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/req
      -- 
    req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(531), ack => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_0); -- 
    concat_cp_element_group_531: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_531"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(514) & concat_CP_34_elements(533);
      gj_concat_cp_element_group_531 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(531), clk => clk, reset => reset); --
    end block;
    -- CP-element group 532:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: marked-predecessors 
    -- CP-element group 532: 	534 
    -- CP-element group 532: 	545 
    -- CP-element group 532: 	556 
    -- CP-element group 532: 	568 
    -- CP-element group 532: 	579 
    -- CP-element group 532: 	615 
    -- CP-element group 532: 	619 
    -- CP-element group 532: 	623 
    -- CP-element group 532: 	627 
    -- CP-element group 532: 	631 
    -- CP-element group 532: 	635 
    -- CP-element group 532: 	647 
    -- CP-element group 532: 	651 
    -- CP-element group 532: 	675 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	534 
    -- CP-element group 532:  members (3) 
      -- CP-element group 532: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_update_start_
      -- CP-element group 532: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/$entry
      -- CP-element group 532: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/req
      -- 
    req_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(532), ack => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_1); -- 
    concat_cp_element_group_532: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_532"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= concat_CP_34_elements(534) & concat_CP_34_elements(545) & concat_CP_34_elements(556) & concat_CP_34_elements(568) & concat_CP_34_elements(579) & concat_CP_34_elements(615) & concat_CP_34_elements(619) & concat_CP_34_elements(623) & concat_CP_34_elements(627) & concat_CP_34_elements(631) & concat_CP_34_elements(635) & concat_CP_34_elements(647) & concat_CP_34_elements(651) & concat_CP_34_elements(675);
      gj_concat_cp_element_group_532 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(532), clk => clk, reset => reset); --
    end block;
    -- CP-element group 533:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	531 
    -- CP-element group 533: successors 
    -- CP-element group 533: marked-successors 
    -- CP-element group 533: 	504 
    -- CP-element group 533: 	512 
    -- CP-element group 533: 	531 
    -- CP-element group 533:  members (3) 
      -- CP-element group 533: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_sample_completed_
      -- CP-element group 533: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/$exit
      -- CP-element group 533: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/ack
      -- 
    ack_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_0, ack => concat_CP_34_elements(533)); -- 
    -- CP-element group 534:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	532 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	543 
    -- CP-element group 534: 	554 
    -- CP-element group 534: 	566 
    -- CP-element group 534: 	577 
    -- CP-element group 534: 	613 
    -- CP-element group 534: 	617 
    -- CP-element group 534: 	621 
    -- CP-element group 534: 	625 
    -- CP-element group 534: 	629 
    -- CP-element group 534: 	633 
    -- CP-element group 534: 	645 
    -- CP-element group 534: 	649 
    -- CP-element group 534: 	673 
    -- CP-element group 534: marked-successors 
    -- CP-element group 534: 	532 
    -- CP-element group 534:  members (3) 
      -- CP-element group 534: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_update_completed_
      -- CP-element group 534: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/$exit
      -- CP-element group 534: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/ack
      -- 
    ack_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_1, ack => concat_CP_34_elements(534)); -- 
    -- CP-element group 535:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	506 
    -- CP-element group 535: 	514 
    -- CP-element group 535: marked-predecessors 
    -- CP-element group 535: 	537 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	537 
    -- CP-element group 535:  members (3) 
      -- CP-element group 535: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/req
      -- 
    req_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(535), ack => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_0); -- 
    concat_cp_element_group_535: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_535"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(514) & concat_CP_34_elements(537);
      gj_concat_cp_element_group_535 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(535), clk => clk, reset => reset); --
    end block;
    -- CP-element group 536:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: marked-predecessors 
    -- CP-element group 536: 	538 
    -- CP-element group 536: 	615 
    -- CP-element group 536: 	619 
    -- CP-element group 536: 	623 
    -- CP-element group 536: 	627 
    -- CP-element group 536: 	631 
    -- CP-element group 536: 	635 
    -- CP-element group 536: 	647 
    -- CP-element group 536: 	651 
    -- CP-element group 536: 	675 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	538 
    -- CP-element group 536:  members (3) 
      -- CP-element group 536: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_update_start_
      -- CP-element group 536: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/req
      -- 
    req_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(536), ack => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_1); -- 
    concat_cp_element_group_536: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_536"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= concat_CP_34_elements(538) & concat_CP_34_elements(615) & concat_CP_34_elements(619) & concat_CP_34_elements(623) & concat_CP_34_elements(627) & concat_CP_34_elements(631) & concat_CP_34_elements(635) & concat_CP_34_elements(647) & concat_CP_34_elements(651) & concat_CP_34_elements(675);
      gj_concat_cp_element_group_536 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(536), clk => clk, reset => reset); --
    end block;
    -- CP-element group 537:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	535 
    -- CP-element group 537: successors 
    -- CP-element group 537: marked-successors 
    -- CP-element group 537: 	504 
    -- CP-element group 537: 	512 
    -- CP-element group 537: 	535 
    -- CP-element group 537:  members (3) 
      -- CP-element group 537: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_sample_completed_
      -- CP-element group 537: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/$exit
      -- CP-element group 537: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/ack
      -- 
    ack_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_0, ack => concat_CP_34_elements(537)); -- 
    -- CP-element group 538:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	536 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	613 
    -- CP-element group 538: 	617 
    -- CP-element group 538: 	621 
    -- CP-element group 538: 	625 
    -- CP-element group 538: 	629 
    -- CP-element group 538: 	633 
    -- CP-element group 538: 	645 
    -- CP-element group 538: 	649 
    -- CP-element group 538: 	673 
    -- CP-element group 538: marked-successors 
    -- CP-element group 538: 	536 
    -- CP-element group 538:  members (3) 
      -- CP-element group 538: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_update_completed_
      -- CP-element group 538: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/$exit
      -- CP-element group 538: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/ack
      -- 
    ack_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 538_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_1, ack => concat_CP_34_elements(538)); -- 
    -- CP-element group 539:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	367 
    -- CP-element group 539: marked-predecessors 
    -- CP-element group 539: 	541 
    -- CP-element group 539: successors 
    -- CP-element group 539: 	541 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_sample_start_
      -- CP-element group 539: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/$entry
      -- CP-element group 539: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/req
      -- 
    req_2301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(539), ack => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_0); -- 
    concat_cp_element_group_539: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_539"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(367) & concat_CP_34_elements(541);
      gj_concat_cp_element_group_539 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(539), clk => clk, reset => reset); --
    end block;
    -- CP-element group 540:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: marked-predecessors 
    -- CP-element group 540: 	542 
    -- CP-element group 540: 	545 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	542 
    -- CP-element group 540:  members (3) 
      -- CP-element group 540: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_update_start_
      -- CP-element group 540: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/$entry
      -- CP-element group 540: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/req
      -- 
    req_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(540), ack => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_1); -- 
    concat_cp_element_group_540: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_540"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(542) & concat_CP_34_elements(545);
      gj_concat_cp_element_group_540 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(540), clk => clk, reset => reset); --
    end block;
    -- CP-element group 541:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	539 
    -- CP-element group 541: successors 
    -- CP-element group 541: marked-successors 
    -- CP-element group 541: 	363 
    -- CP-element group 541: 	539 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_sample_completed_
      -- CP-element group 541: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/$exit
      -- CP-element group 541: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/ack
      -- 
    ack_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_0, ack => concat_CP_34_elements(541)); -- 
    -- CP-element group 542:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	540 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	543 
    -- CP-element group 542: marked-successors 
    -- CP-element group 542: 	540 
    -- CP-element group 542:  members (3) 
      -- CP-element group 542: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_update_completed_
      -- CP-element group 542: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/$exit
      -- CP-element group 542: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/ack
      -- 
    ack_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 542_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_1, ack => concat_CP_34_elements(542)); -- 
    -- CP-element group 543:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	526 
    -- CP-element group 543: 	534 
    -- CP-element group 543: 	542 
    -- CP-element group 543: marked-predecessors 
    -- CP-element group 543: 	545 
    -- CP-element group 543: successors 
    -- CP-element group 543: 	545 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_sample_start_
      -- CP-element group 543: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/$entry
      -- CP-element group 543: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/rr
      -- 
    rr_2315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(543), ack => type_cast_1073_inst_req_0); -- 
    concat_cp_element_group_543: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_543"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(542) & concat_CP_34_elements(545);
      gj_concat_cp_element_group_543 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(543), clk => clk, reset => reset); --
    end block;
    -- CP-element group 544:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: marked-predecessors 
    -- CP-element group 544: 	546 
    -- CP-element group 544: 	550 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	546 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_update_start_
      -- CP-element group 544: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/$entry
      -- CP-element group 544: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/cr
      -- 
    cr_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(544), ack => type_cast_1073_inst_req_1); -- 
    concat_cp_element_group_544: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_544"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(546) & concat_CP_34_elements(550);
      gj_concat_cp_element_group_544 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(544), clk => clk, reset => reset); --
    end block;
    -- CP-element group 545:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	543 
    -- CP-element group 545: successors 
    -- CP-element group 545: marked-successors 
    -- CP-element group 545: 	524 
    -- CP-element group 545: 	532 
    -- CP-element group 545: 	540 
    -- CP-element group 545: 	543 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_sample_completed_
      -- CP-element group 545: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/$exit
      -- CP-element group 545: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/ra
      -- 
    ra_2316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 545_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_0, ack => concat_CP_34_elements(545)); -- 
    -- CP-element group 546:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	544 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	550 
    -- CP-element group 546: marked-successors 
    -- CP-element group 546: 	544 
    -- CP-element group 546:  members (16) 
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_update_completed_
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/$exit
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/ca
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resized_1
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scaled_1
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_computed_1
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/$entry
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/$exit
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/index_resize_req
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/index_resize_ack
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/$entry
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/$exit
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/scale_rename_req
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/scale_rename_ack
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/$entry
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/req
      -- 
    ca_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_1, ack => concat_CP_34_elements(546)); -- 
    req_2346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(546), ack => array_obj_ref_1079_index_offset_req_0); -- 
    -- CP-element group 547:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	551 
    -- CP-element group 547: marked-predecessors 
    -- CP-element group 547: 	552 
    -- CP-element group 547: successors 
    -- CP-element group 547: 	552 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_sample_start_
      -- CP-element group 547: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/$entry
      -- CP-element group 547: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/req
      -- 
    req_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(547), ack => addr_of_1080_final_reg_req_0); -- 
    concat_cp_element_group_547: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_547"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(551) & concat_CP_34_elements(552);
      gj_concat_cp_element_group_547 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(547), clk => clk, reset => reset); --
    end block;
    -- CP-element group 548:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	316 
    -- CP-element group 548: marked-predecessors 
    -- CP-element group 548: 	553 
    -- CP-element group 548: 	560 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	553 
    -- CP-element group 548:  members (3) 
      -- CP-element group 548: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_update_start_
      -- CP-element group 548: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/$entry
      -- CP-element group 548: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/req
      -- 
    req_2366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(548), ack => addr_of_1080_final_reg_req_1); -- 
    concat_cp_element_group_548: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_548"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(553) & concat_CP_34_elements(560);
      gj_concat_cp_element_group_548 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(548), clk => clk, reset => reset); --
    end block;
    -- CP-element group 549:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	316 
    -- CP-element group 549: marked-predecessors 
    -- CP-element group 549: 	551 
    -- CP-element group 549: 	552 
    -- CP-element group 549: successors 
    -- CP-element group 549: 	551 
    -- CP-element group 549:  members (3) 
      -- CP-element group 549: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_update_start
      -- CP-element group 549: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/$entry
      -- CP-element group 549: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/req
      -- 
    req_2351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(549), ack => array_obj_ref_1079_index_offset_req_1); -- 
    concat_cp_element_group_549: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_549"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(551) & concat_CP_34_elements(552);
      gj_concat_cp_element_group_549 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(549), clk => clk, reset => reset); --
    end block;
    -- CP-element group 550:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	546 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	691 
    -- CP-element group 550: marked-successors 
    -- CP-element group 550: 	544 
    -- CP-element group 550:  members (3) 
      -- CP-element group 550: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_sample_complete
      -- CP-element group 550: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/$exit
      -- CP-element group 550: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/ack
      -- 
    ack_2347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_index_offset_ack_0, ack => concat_CP_34_elements(550)); -- 
    -- CP-element group 551:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	549 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	547 
    -- CP-element group 551: marked-successors 
    -- CP-element group 551: 	549 
    -- CP-element group 551:  members (8) 
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_root_address_calculated
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_offset_calculated
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/$exit
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/ack
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/$entry
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/$exit
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/sum_rename_req
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/sum_rename_ack
      -- 
    ack_2352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 551_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_index_offset_ack_1, ack => concat_CP_34_elements(551)); -- 
    -- CP-element group 552:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	547 
    -- CP-element group 552: successors 
    -- CP-element group 552: marked-successors 
    -- CP-element group 552: 	547 
    -- CP-element group 552: 	549 
    -- CP-element group 552:  members (3) 
      -- CP-element group 552: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_sample_completed_
      -- CP-element group 552: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/$exit
      -- CP-element group 552: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/ack
      -- 
    ack_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1080_final_reg_ack_0, ack => concat_CP_34_elements(552)); -- 
    -- CP-element group 553:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	548 
    -- CP-element group 553: successors 
    -- CP-element group 553: 	558 
    -- CP-element group 553: marked-successors 
    -- CP-element group 553: 	548 
    -- CP-element group 553:  members (19) 
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_update_completed_
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/$exit
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/ack
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_address_calculated
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_address_calculated
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_root_address_calculated
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_address_resized
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/$entry
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/$exit
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/base_resize_req
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/base_resize_ack
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/$entry
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/$exit
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/sum_rename_req
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/sum_rename_ack
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/$entry
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/$exit
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/root_register_req
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/root_register_ack
      -- 
    ack_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1080_final_reg_ack_1, ack => concat_CP_34_elements(553)); -- 
    -- CP-element group 554:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	526 
    -- CP-element group 554: 	534 
    -- CP-element group 554: marked-predecessors 
    -- CP-element group 554: 	556 
    -- CP-element group 554: successors 
    -- CP-element group 554: 	556 
    -- CP-element group 554:  members (3) 
      -- CP-element group 554: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_sample_start_
      -- CP-element group 554: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/$entry
      -- CP-element group 554: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/req
      -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(554), ack => W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_req_0); -- 
    concat_cp_element_group_554: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_554"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(556);
      gj_concat_cp_element_group_554 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(554), clk => clk, reset => reset); --
    end block;
    -- CP-element group 555:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: marked-predecessors 
    -- CP-element group 555: 	557 
    -- CP-element group 555: 	560 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	557 
    -- CP-element group 555:  members (3) 
      -- CP-element group 555: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_update_start_
      -- CP-element group 555: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/$entry
      -- CP-element group 555: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/req
      -- 
    req_2380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(555), ack => W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_req_1); -- 
    concat_cp_element_group_555: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_555"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(557) & concat_CP_34_elements(560);
      gj_concat_cp_element_group_555 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(555), clk => clk, reset => reset); --
    end block;
    -- CP-element group 556:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	554 
    -- CP-element group 556: successors 
    -- CP-element group 556: marked-successors 
    -- CP-element group 556: 	524 
    -- CP-element group 556: 	532 
    -- CP-element group 556: 	554 
    -- CP-element group 556:  members (3) 
      -- CP-element group 556: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_sample_completed_
      -- CP-element group 556: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/$exit
      -- CP-element group 556: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/ack
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_ack_0, ack => concat_CP_34_elements(556)); -- 
    -- CP-element group 557:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	555 
    -- CP-element group 557: successors 
    -- CP-element group 557: 	558 
    -- CP-element group 557: marked-successors 
    -- CP-element group 557: 	555 
    -- CP-element group 557:  members (3) 
      -- CP-element group 557: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_update_completed_
      -- CP-element group 557: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/$exit
      -- CP-element group 557: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/ack
      -- 
    ack_2381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_ack_1, ack => concat_CP_34_elements(557)); -- 
    -- CP-element group 558:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	553 
    -- CP-element group 558: 	557 
    -- CP-element group 558: marked-predecessors 
    -- CP-element group 558: 	560 
    -- CP-element group 558: successors 
    -- CP-element group 558: 	560 
    -- CP-element group 558:  members (5) 
      -- CP-element group 558: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_sample_start_
      -- CP-element group 558: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/rr
      -- 
    rr_2414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => ptr_deref_1088_load_0_req_0); -- 
    concat_cp_element_group_558: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_558"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(553) & concat_CP_34_elements(557) & concat_CP_34_elements(560);
      gj_concat_cp_element_group_558 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(558), clk => clk, reset => reset); --
    end block;
    -- CP-element group 559:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: marked-predecessors 
    -- CP-element group 559: 	561 
    -- CP-element group 559: 	587 
    -- CP-element group 559: successors 
    -- CP-element group 559: 	561 
    -- CP-element group 559:  members (5) 
      -- CP-element group 559: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_update_start_
      -- CP-element group 559: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/$entry
      -- CP-element group 559: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/$entry
      -- CP-element group 559: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/cr
      -- 
    cr_2425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(559), ack => ptr_deref_1088_load_0_req_1); -- 
    concat_cp_element_group_559: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_559"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(561) & concat_CP_34_elements(587);
      gj_concat_cp_element_group_559 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(559), clk => clk, reset => reset); --
    end block;
    -- CP-element group 560:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	558 
    -- CP-element group 560: successors 
    -- CP-element group 560: marked-successors 
    -- CP-element group 560: 	548 
    -- CP-element group 560: 	555 
    -- CP-element group 560: 	558 
    -- CP-element group 560:  members (5) 
      -- CP-element group 560: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_sample_completed_
      -- CP-element group 560: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/$exit
      -- CP-element group 560: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/$exit
      -- CP-element group 560: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/$exit
      -- CP-element group 560: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/ra
      -- 
    ra_2415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 560_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_load_0_ack_0, ack => concat_CP_34_elements(560)); -- 
    -- CP-element group 561:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	559 
    -- CP-element group 561: successors 
    -- CP-element group 561: 	585 
    -- CP-element group 561: marked-successors 
    -- CP-element group 561: 	559 
    -- CP-element group 561:  members (9) 
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_update_completed_
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/$exit
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/$exit
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/$exit
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/ca
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/$entry
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/$exit
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/merge_req
      -- CP-element group 561: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/merge_ack
      -- 
    ca_2426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 561_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_load_0_ack_1, ack => concat_CP_34_elements(561)); -- 
    -- CP-element group 562:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	428 
    -- CP-element group 562: 	490 
    -- CP-element group 562: 	494 
    -- CP-element group 562: marked-predecessors 
    -- CP-element group 562: 	564 
    -- CP-element group 562: successors 
    -- CP-element group 562: 	564 
    -- CP-element group 562:  members (3) 
      -- CP-element group 562: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/req
      -- 
    req_2439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => W_add_outx_x0_1032_delayed_2_0_1090_inst_req_0); -- 
    concat_cp_element_group_562: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_562"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(490) & concat_CP_34_elements(494) & concat_CP_34_elements(564);
      gj_concat_cp_element_group_562 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(562), clk => clk, reset => reset); --
    end block;
    -- CP-element group 563:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: marked-predecessors 
    -- CP-element group 563: 	565 
    -- CP-element group 563: 	568 
    -- CP-element group 563: successors 
    -- CP-element group 563: 	565 
    -- CP-element group 563:  members (3) 
      -- CP-element group 563: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_update_start_
      -- CP-element group 563: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/$entry
      -- CP-element group 563: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/req
      -- 
    req_2444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(563), ack => W_add_outx_x0_1032_delayed_2_0_1090_inst_req_1); -- 
    concat_cp_element_group_563: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_563"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(565) & concat_CP_34_elements(568);
      gj_concat_cp_element_group_563 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(563), clk => clk, reset => reset); --
    end block;
    -- CP-element group 564:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	562 
    -- CP-element group 564: successors 
    -- CP-element group 564: marked-successors 
    -- CP-element group 564: 	426 
    -- CP-element group 564: 	488 
    -- CP-element group 564: 	492 
    -- CP-element group 564: 	562 
    -- CP-element group 564:  members (3) 
      -- CP-element group 564: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_sample_completed_
      -- CP-element group 564: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/$exit
      -- CP-element group 564: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/ack
      -- 
    ack_2440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 564_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_0, ack => concat_CP_34_elements(564)); -- 
    -- CP-element group 565:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	563 
    -- CP-element group 565: successors 
    -- CP-element group 565: 	566 
    -- CP-element group 565: marked-successors 
    -- CP-element group 565: 	563 
    -- CP-element group 565:  members (3) 
      -- CP-element group 565: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_update_completed_
      -- CP-element group 565: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/$exit
      -- CP-element group 565: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/ack
      -- 
    ack_2445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_1, ack => concat_CP_34_elements(565)); -- 
    -- CP-element group 566:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	526 
    -- CP-element group 566: 	534 
    -- CP-element group 566: 	565 
    -- CP-element group 566: marked-predecessors 
    -- CP-element group 566: 	568 
    -- CP-element group 566: successors 
    -- CP-element group 566: 	568 
    -- CP-element group 566:  members (3) 
      -- CP-element group 566: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_sample_start_
      -- CP-element group 566: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/$entry
      -- CP-element group 566: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/rr
      -- 
    rr_2453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(566), ack => type_cast_1096_inst_req_0); -- 
    concat_cp_element_group_566: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_566"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(565) & concat_CP_34_elements(568);
      gj_concat_cp_element_group_566 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(566), clk => clk, reset => reset); --
    end block;
    -- CP-element group 567:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: marked-predecessors 
    -- CP-element group 567: 	569 
    -- CP-element group 567: 	573 
    -- CP-element group 567: successors 
    -- CP-element group 567: 	569 
    -- CP-element group 567:  members (3) 
      -- CP-element group 567: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_update_start_
      -- CP-element group 567: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/$entry
      -- CP-element group 567: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/cr
      -- 
    cr_2458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(567), ack => type_cast_1096_inst_req_1); -- 
    concat_cp_element_group_567: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_567"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(569) & concat_CP_34_elements(573);
      gj_concat_cp_element_group_567 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(567), clk => clk, reset => reset); --
    end block;
    -- CP-element group 568:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	566 
    -- CP-element group 568: successors 
    -- CP-element group 568: marked-successors 
    -- CP-element group 568: 	524 
    -- CP-element group 568: 	532 
    -- CP-element group 568: 	563 
    -- CP-element group 568: 	566 
    -- CP-element group 568:  members (3) 
      -- CP-element group 568: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_sample_completed_
      -- CP-element group 568: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/$exit
      -- CP-element group 568: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/ra
      -- 
    ra_2454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 568_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1096_inst_ack_0, ack => concat_CP_34_elements(568)); -- 
    -- CP-element group 569:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	567 
    -- CP-element group 569: successors 
    -- CP-element group 569: 	573 
    -- CP-element group 569: marked-successors 
    -- CP-element group 569: 	567 
    -- CP-element group 569:  members (16) 
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_update_completed_
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/$exit
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/ca
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resized_1
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scaled_1
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_computed_1
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/$entry
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/$exit
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/index_resize_req
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/index_resize_ack
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/$entry
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/$exit
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/scale_rename_req
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/scale_rename_ack
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/$entry
      -- CP-element group 569: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/req
      -- 
    ca_2459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 569_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1096_inst_ack_1, ack => concat_CP_34_elements(569)); -- 
    req_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(569), ack => array_obj_ref_1102_index_offset_req_0); -- 
    -- CP-element group 570:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: 	574 
    -- CP-element group 570: marked-predecessors 
    -- CP-element group 570: 	575 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	575 
    -- CP-element group 570:  members (3) 
      -- CP-element group 570: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_sample_start_
      -- CP-element group 570: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/$entry
      -- CP-element group 570: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/req
      -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(570), ack => addr_of_1103_final_reg_req_0); -- 
    concat_cp_element_group_570: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_570"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(574) & concat_CP_34_elements(575);
      gj_concat_cp_element_group_570 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(570), clk => clk, reset => reset); --
    end block;
    -- CP-element group 571:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	316 
    -- CP-element group 571: marked-predecessors 
    -- CP-element group 571: 	576 
    -- CP-element group 571: 	583 
    -- CP-element group 571: successors 
    -- CP-element group 571: 	576 
    -- CP-element group 571:  members (3) 
      -- CP-element group 571: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_update_start_
      -- CP-element group 571: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/$entry
      -- CP-element group 571: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/req
      -- 
    req_2504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(571), ack => addr_of_1103_final_reg_req_1); -- 
    concat_cp_element_group_571: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_571"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(576) & concat_CP_34_elements(583);
      gj_concat_cp_element_group_571 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(571), clk => clk, reset => reset); --
    end block;
    -- CP-element group 572:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	316 
    -- CP-element group 572: marked-predecessors 
    -- CP-element group 572: 	574 
    -- CP-element group 572: 	575 
    -- CP-element group 572: successors 
    -- CP-element group 572: 	574 
    -- CP-element group 572:  members (3) 
      -- CP-element group 572: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_update_start
      -- CP-element group 572: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/$entry
      -- CP-element group 572: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/req
      -- 
    req_2489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(572), ack => array_obj_ref_1102_index_offset_req_1); -- 
    concat_cp_element_group_572: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_572"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(574) & concat_CP_34_elements(575);
      gj_concat_cp_element_group_572 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(572), clk => clk, reset => reset); --
    end block;
    -- CP-element group 573:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	569 
    -- CP-element group 573: successors 
    -- CP-element group 573: 	691 
    -- CP-element group 573: marked-successors 
    -- CP-element group 573: 	567 
    -- CP-element group 573:  members (3) 
      -- CP-element group 573: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_sample_complete
      -- CP-element group 573: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/$exit
      -- CP-element group 573: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/ack
      -- 
    ack_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 573_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1102_index_offset_ack_0, ack => concat_CP_34_elements(573)); -- 
    -- CP-element group 574:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	572 
    -- CP-element group 574: successors 
    -- CP-element group 574: 	570 
    -- CP-element group 574: marked-successors 
    -- CP-element group 574: 	572 
    -- CP-element group 574:  members (8) 
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_root_address_calculated
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_offset_calculated
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/$exit
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/ack
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/$entry
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/$exit
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/sum_rename_req
      -- CP-element group 574: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/sum_rename_ack
      -- 
    ack_2490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 574_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1102_index_offset_ack_1, ack => concat_CP_34_elements(574)); -- 
    -- CP-element group 575:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	570 
    -- CP-element group 575: successors 
    -- CP-element group 575: marked-successors 
    -- CP-element group 575: 	570 
    -- CP-element group 575: 	572 
    -- CP-element group 575:  members (3) 
      -- CP-element group 575: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_sample_completed_
      -- CP-element group 575: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/$exit
      -- CP-element group 575: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/ack
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 575_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1103_final_reg_ack_0, ack => concat_CP_34_elements(575)); -- 
    -- CP-element group 576:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	571 
    -- CP-element group 576: successors 
    -- CP-element group 576: 	581 
    -- CP-element group 576: marked-successors 
    -- CP-element group 576: 	571 
    -- CP-element group 576:  members (3) 
      -- CP-element group 576: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_update_completed_
      -- CP-element group 576: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/$exit
      -- CP-element group 576: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/ack
      -- 
    ack_2505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 576_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1103_final_reg_ack_1, ack => concat_CP_34_elements(576)); -- 
    -- CP-element group 577:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	526 
    -- CP-element group 577: 	534 
    -- CP-element group 577: marked-predecessors 
    -- CP-element group 577: 	579 
    -- CP-element group 577: successors 
    -- CP-element group 577: 	579 
    -- CP-element group 577:  members (3) 
      -- CP-element group 577: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_sample_start_
      -- CP-element group 577: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/$entry
      -- CP-element group 577: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/req
      -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(577), ack => W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_req_0); -- 
    concat_cp_element_group_577: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_577"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(579);
      gj_concat_cp_element_group_577 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(577), clk => clk, reset => reset); --
    end block;
    -- CP-element group 578:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: marked-predecessors 
    -- CP-element group 578: 	580 
    -- CP-element group 578: successors 
    -- CP-element group 578: 	580 
    -- CP-element group 578:  members (3) 
      -- CP-element group 578: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_update_start_
      -- CP-element group 578: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/$entry
      -- CP-element group 578: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/req
      -- 
    req_2518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(578), ack => W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_req_1); -- 
    concat_cp_element_group_578: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_578"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(580);
      gj_concat_cp_element_group_578 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(578), clk => clk, reset => reset); --
    end block;
    -- CP-element group 579:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	577 
    -- CP-element group 579: successors 
    -- CP-element group 579: marked-successors 
    -- CP-element group 579: 	524 
    -- CP-element group 579: 	532 
    -- CP-element group 579: 	577 
    -- CP-element group 579:  members (3) 
      -- CP-element group 579: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_sample_completed_
      -- CP-element group 579: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/$exit
      -- CP-element group 579: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/ack
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 579_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_ack_0, ack => concat_CP_34_elements(579)); -- 
    -- CP-element group 580:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	578 
    -- CP-element group 580: successors 
    -- CP-element group 580: 	691 
    -- CP-element group 580: marked-successors 
    -- CP-element group 580: 	578 
    -- CP-element group 580:  members (3) 
      -- CP-element group 580: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_update_completed_
      -- CP-element group 580: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/$exit
      -- CP-element group 580: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/ack
      -- 
    ack_2519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 580_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_ack_1, ack => concat_CP_34_elements(580)); -- 
    -- CP-element group 581:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	576 
    -- CP-element group 581: marked-predecessors 
    -- CP-element group 581: 	583 
    -- CP-element group 581: successors 
    -- CP-element group 581: 	583 
    -- CP-element group 581:  members (3) 
      -- CP-element group 581: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_sample_start_
      -- CP-element group 581: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/$entry
      -- CP-element group 581: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/req
      -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(581), ack => W_arrayidx273_1043_delayed_6_0_1108_inst_req_0); -- 
    concat_cp_element_group_581: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_581"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(576) & concat_CP_34_elements(583);
      gj_concat_cp_element_group_581 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(581), clk => clk, reset => reset); --
    end block;
    -- CP-element group 582:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: marked-predecessors 
    -- CP-element group 582: 	584 
    -- CP-element group 582: 	587 
    -- CP-element group 582: successors 
    -- CP-element group 582: 	584 
    -- CP-element group 582:  members (3) 
      -- CP-element group 582: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_update_start_
      -- CP-element group 582: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/$entry
      -- CP-element group 582: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/req
      -- 
    req_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(582), ack => W_arrayidx273_1043_delayed_6_0_1108_inst_req_1); -- 
    concat_cp_element_group_582: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_582"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(584) & concat_CP_34_elements(587);
      gj_concat_cp_element_group_582 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(582), clk => clk, reset => reset); --
    end block;
    -- CP-element group 583:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	581 
    -- CP-element group 583: successors 
    -- CP-element group 583: marked-successors 
    -- CP-element group 583: 	571 
    -- CP-element group 583: 	581 
    -- CP-element group 583:  members (3) 
      -- CP-element group 583: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_sample_completed_
      -- CP-element group 583: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/$exit
      -- CP-element group 583: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/ack
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx273_1043_delayed_6_0_1108_inst_ack_0, ack => concat_CP_34_elements(583)); -- 
    -- CP-element group 584:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	582 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	585 
    -- CP-element group 584: marked-successors 
    -- CP-element group 584: 	582 
    -- CP-element group 584:  members (19) 
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_update_completed_
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/$exit
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/ack
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_address_calculated
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_address_calculated
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_root_address_calculated
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_address_resized
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/$entry
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/$exit
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/base_resize_req
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/base_resize_ack
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/$entry
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/$exit
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/sum_rename_req
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/sum_rename_ack
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/$entry
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/$exit
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/root_register_req
      -- CP-element group 584: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/root_register_ack
      -- 
    ack_2533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 584_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx273_1043_delayed_6_0_1108_inst_ack_1, ack => concat_CP_34_elements(584)); -- 
    -- CP-element group 585:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	561 
    -- CP-element group 585: 	584 
    -- CP-element group 585: 	690 
    -- CP-element group 585: marked-predecessors 
    -- CP-element group 585: 	587 
    -- CP-element group 585: successors 
    -- CP-element group 585: 	587 
    -- CP-element group 585:  members (9) 
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_sample_start_
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/$entry
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/$entry
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/$exit
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/split_req
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/split_ack
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/$entry
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/$entry
      -- CP-element group 585: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/rr
      -- 
    rr_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(585), ack => ptr_deref_1113_store_0_req_0); -- 
    concat_cp_element_group_585: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_585"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(561) & concat_CP_34_elements(584) & concat_CP_34_elements(690) & concat_CP_34_elements(587);
      gj_concat_cp_element_group_585 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(585), clk => clk, reset => reset); --
    end block;
    -- CP-element group 586:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: marked-predecessors 
    -- CP-element group 586: 	588 
    -- CP-element group 586: successors 
    -- CP-element group 586: 	588 
    -- CP-element group 586:  members (5) 
      -- CP-element group 586: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_update_start_
      -- CP-element group 586: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/$entry
      -- CP-element group 586: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/$entry
      -- CP-element group 586: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/$entry
      -- CP-element group 586: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/cr
      -- 
    cr_2582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(586), ack => ptr_deref_1113_store_0_req_1); -- 
    concat_cp_element_group_586: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_586"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(588);
      gj_concat_cp_element_group_586 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(586), clk => clk, reset => reset); --
    end block;
    -- CP-element group 587:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	585 
    -- CP-element group 587: successors 
    -- CP-element group 587: 	691 
    -- CP-element group 587: marked-successors 
    -- CP-element group 587: 	475 
    -- CP-element group 587: 	559 
    -- CP-element group 587: 	582 
    -- CP-element group 587: 	585 
    -- CP-element group 587:  members (6) 
      -- CP-element group 587: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_sample_completed_
      -- CP-element group 587: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/$exit
      -- CP-element group 587: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/$exit
      -- CP-element group 587: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/$exit
      -- CP-element group 587: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/ra
      -- CP-element group 587: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ring_reenable_memory_space_2
      -- 
    ra_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 587_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_store_0_ack_0, ack => concat_CP_34_elements(587)); -- 
    -- CP-element group 588:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	586 
    -- CP-element group 588: successors 
    -- CP-element group 588: 	691 
    -- CP-element group 588: marked-successors 
    -- CP-element group 588: 	586 
    -- CP-element group 588:  members (5) 
      -- CP-element group 588: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_update_completed_
      -- CP-element group 588: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/$exit
      -- CP-element group 588: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/$exit
      -- CP-element group 588: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/$exit
      -- CP-element group 588: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/ca
      -- 
    ca_2583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 588_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_store_0_ack_1, ack => concat_CP_34_elements(588)); -- 
    -- CP-element group 589:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	409 
    -- CP-element group 589: marked-predecessors 
    -- CP-element group 589: 	591 
    -- CP-element group 589: successors 
    -- CP-element group 589: 	591 
    -- CP-element group 589:  members (3) 
      -- CP-element group 589: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_sample_start_
      -- CP-element group 589: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/$entry
      -- CP-element group 589: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/req
      -- 
    req_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(589), ack => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_0); -- 
    concat_cp_element_group_589: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_589"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(409) & concat_CP_34_elements(591);
      gj_concat_cp_element_group_589 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(589), clk => clk, reset => reset); --
    end block;
    -- CP-element group 590:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: marked-predecessors 
    -- CP-element group 590: 	592 
    -- CP-element group 590: 	615 
    -- CP-element group 590: 	675 
    -- CP-element group 590: successors 
    -- CP-element group 590: 	592 
    -- CP-element group 590:  members (3) 
      -- CP-element group 590: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_update_start_
      -- CP-element group 590: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/$entry
      -- CP-element group 590: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/req
      -- 
    req_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(590), ack => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_1); -- 
    concat_cp_element_group_590: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_590"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(592) & concat_CP_34_elements(615) & concat_CP_34_elements(675);
      gj_concat_cp_element_group_590 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(590), clk => clk, reset => reset); --
    end block;
    -- CP-element group 591:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	589 
    -- CP-element group 591: successors 
    -- CP-element group 591: marked-successors 
    -- CP-element group 591: 	405 
    -- CP-element group 591: 	589 
    -- CP-element group 591:  members (3) 
      -- CP-element group 591: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_sample_completed_
      -- CP-element group 591: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/$exit
      -- CP-element group 591: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/ack
      -- 
    ack_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 591_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_0, ack => concat_CP_34_elements(591)); -- 
    -- CP-element group 592:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	590 
    -- CP-element group 592: successors 
    -- CP-element group 592: 	613 
    -- CP-element group 592: 	673 
    -- CP-element group 592: marked-successors 
    -- CP-element group 592: 	590 
    -- CP-element group 592:  members (3) 
      -- CP-element group 592: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_update_completed_
      -- CP-element group 592: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/$exit
      -- CP-element group 592: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/ack
      -- 
    ack_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 592_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_1, ack => concat_CP_34_elements(592)); -- 
    -- CP-element group 593:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	367 
    -- CP-element group 593: marked-predecessors 
    -- CP-element group 593: 	595 
    -- CP-element group 593: successors 
    -- CP-element group 593: 	595 
    -- CP-element group 593:  members (3) 
      -- CP-element group 593: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_sample_start_
      -- CP-element group 593: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/$entry
      -- CP-element group 593: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/req
      -- 
    req_2605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(593), ack => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_0); -- 
    concat_cp_element_group_593: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_593"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(367) & concat_CP_34_elements(595);
      gj_concat_cp_element_group_593 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(593), clk => clk, reset => reset); --
    end block;
    -- CP-element group 594:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: marked-predecessors 
    -- CP-element group 594: 	596 
    -- CP-element group 594: 	631 
    -- CP-element group 594: 	635 
    -- CP-element group 594: successors 
    -- CP-element group 594: 	596 
    -- CP-element group 594:  members (3) 
      -- CP-element group 594: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_update_start_
      -- CP-element group 594: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/$entry
      -- CP-element group 594: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/req
      -- 
    req_2610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(594), ack => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_1); -- 
    concat_cp_element_group_594: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_594"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(596) & concat_CP_34_elements(631) & concat_CP_34_elements(635);
      gj_concat_cp_element_group_594 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(594), clk => clk, reset => reset); --
    end block;
    -- CP-element group 595:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	593 
    -- CP-element group 595: successors 
    -- CP-element group 595: marked-successors 
    -- CP-element group 595: 	363 
    -- CP-element group 595: 	593 
    -- CP-element group 595:  members (3) 
      -- CP-element group 595: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_sample_completed_
      -- CP-element group 595: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/$exit
      -- CP-element group 595: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/ack
      -- 
    ack_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 595_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_0, ack => concat_CP_34_elements(595)); -- 
    -- CP-element group 596:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	594 
    -- CP-element group 596: successors 
    -- CP-element group 596: 	629 
    -- CP-element group 596: 	633 
    -- CP-element group 596: marked-successors 
    -- CP-element group 596: 	594 
    -- CP-element group 596:  members (3) 
      -- CP-element group 596: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_update_completed_
      -- CP-element group 596: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/$exit
      -- CP-element group 596: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/ack
      -- 
    ack_2611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 596_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_1, ack => concat_CP_34_elements(596)); -- 
    -- CP-element group 597:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	428 
    -- CP-element group 597: 	490 
    -- CP-element group 597: 	494 
    -- CP-element group 597: marked-predecessors 
    -- CP-element group 597: 	599 
    -- CP-element group 597: successors 
    -- CP-element group 597: 	599 
    -- CP-element group 597:  members (3) 
      -- CP-element group 597: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_sample_start_
      -- CP-element group 597: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/$entry
      -- CP-element group 597: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/req
      -- 
    req_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(597), ack => W_add_outx_x0_1063_delayed_2_0_1136_inst_req_0); -- 
    concat_cp_element_group_597: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_597"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(490) & concat_CP_34_elements(494) & concat_CP_34_elements(599);
      gj_concat_cp_element_group_597 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(597), clk => clk, reset => reset); --
    end block;
    -- CP-element group 598:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: marked-predecessors 
    -- CP-element group 598: 	600 
    -- CP-element group 598: 	647 
    -- CP-element group 598: 	651 
    -- CP-element group 598: successors 
    -- CP-element group 598: 	600 
    -- CP-element group 598:  members (3) 
      -- CP-element group 598: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_update_start_
      -- CP-element group 598: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/$entry
      -- CP-element group 598: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/req
      -- 
    req_2624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(598), ack => W_add_outx_x0_1063_delayed_2_0_1136_inst_req_1); -- 
    concat_cp_element_group_598: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_598"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(600) & concat_CP_34_elements(647) & concat_CP_34_elements(651);
      gj_concat_cp_element_group_598 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(598), clk => clk, reset => reset); --
    end block;
    -- CP-element group 599:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	597 
    -- CP-element group 599: successors 
    -- CP-element group 599: marked-successors 
    -- CP-element group 599: 	426 
    -- CP-element group 599: 	488 
    -- CP-element group 599: 	492 
    -- CP-element group 599: 	597 
    -- CP-element group 599:  members (3) 
      -- CP-element group 599: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_sample_completed_
      -- CP-element group 599: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/$exit
      -- CP-element group 599: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/ack
      -- 
    ack_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 599_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_0, ack => concat_CP_34_elements(599)); -- 
    -- CP-element group 600:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	598 
    -- CP-element group 600: successors 
    -- CP-element group 600: 	645 
    -- CP-element group 600: 	649 
    -- CP-element group 600: marked-successors 
    -- CP-element group 600: 	598 
    -- CP-element group 600:  members (3) 
      -- CP-element group 600: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_update_completed_
      -- CP-element group 600: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/$exit
      -- CP-element group 600: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/ack
      -- 
    ack_2625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 600_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_1, ack => concat_CP_34_elements(600)); -- 
    -- CP-element group 601:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	428 
    -- CP-element group 601: 	490 
    -- CP-element group 601: 	494 
    -- CP-element group 601: marked-predecessors 
    -- CP-element group 601: 	603 
    -- CP-element group 601: successors 
    -- CP-element group 601: 	603 
    -- CP-element group 601:  members (3) 
      -- CP-element group 601: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_sample_start_
      -- CP-element group 601: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/$entry
      -- CP-element group 601: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/rr
      -- 
    rr_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(601), ack => type_cast_1156_inst_req_0); -- 
    concat_cp_element_group_601: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_601"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(490) & concat_CP_34_elements(494) & concat_CP_34_elements(603);
      gj_concat_cp_element_group_601 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(601), clk => clk, reset => reset); --
    end block;
    -- CP-element group 602:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: marked-predecessors 
    -- CP-element group 602: 	604 
    -- CP-element group 602: 	647 
    -- CP-element group 602: 	651 
    -- CP-element group 602: successors 
    -- CP-element group 602: 	604 
    -- CP-element group 602:  members (3) 
      -- CP-element group 602: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_update_start_
      -- CP-element group 602: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/$entry
      -- CP-element group 602: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/cr
      -- 
    cr_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(602), ack => type_cast_1156_inst_req_1); -- 
    concat_cp_element_group_602: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_602"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(604) & concat_CP_34_elements(647) & concat_CP_34_elements(651);
      gj_concat_cp_element_group_602 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(602), clk => clk, reset => reset); --
    end block;
    -- CP-element group 603:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	601 
    -- CP-element group 603: successors 
    -- CP-element group 603: marked-successors 
    -- CP-element group 603: 	426 
    -- CP-element group 603: 	488 
    -- CP-element group 603: 	492 
    -- CP-element group 603: 	601 
    -- CP-element group 603:  members (3) 
      -- CP-element group 603: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_sample_completed_
      -- CP-element group 603: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/$exit
      -- CP-element group 603: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/ra
      -- 
    ra_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 603_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_0, ack => concat_CP_34_elements(603)); -- 
    -- CP-element group 604:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	602 
    -- CP-element group 604: successors 
    -- CP-element group 604: 	645 
    -- CP-element group 604: 	649 
    -- CP-element group 604: marked-successors 
    -- CP-element group 604: 	602 
    -- CP-element group 604:  members (3) 
      -- CP-element group 604: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_update_completed_
      -- CP-element group 604: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/$exit
      -- CP-element group 604: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/ca
      -- 
    ca_2639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 604_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_1, ack => concat_CP_34_elements(604)); -- 
    -- CP-element group 605:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	367 
    -- CP-element group 605: marked-predecessors 
    -- CP-element group 605: 	607 
    -- CP-element group 605: successors 
    -- CP-element group 605: 	607 
    -- CP-element group 605:  members (3) 
      -- CP-element group 605: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/$entry
      -- CP-element group 605: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/rr
      -- CP-element group 605: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_sample_start_
      -- 
    rr_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(605), ack => type_cast_1171_inst_req_0); -- 
    concat_cp_element_group_605: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_605"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(367) & concat_CP_34_elements(607);
      gj_concat_cp_element_group_605 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(605), clk => clk, reset => reset); --
    end block;
    -- CP-element group 606:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: marked-predecessors 
    -- CP-element group 606: 	608 
    -- CP-element group 606: 	631 
    -- CP-element group 606: 	635 
    -- CP-element group 606: successors 
    -- CP-element group 606: 	608 
    -- CP-element group 606:  members (3) 
      -- CP-element group 606: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/$entry
      -- CP-element group 606: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/cr
      -- CP-element group 606: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_update_start_
      -- 
    cr_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(606), ack => type_cast_1171_inst_req_1); -- 
    concat_cp_element_group_606: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_606"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(608) & concat_CP_34_elements(631) & concat_CP_34_elements(635);
      gj_concat_cp_element_group_606 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(606), clk => clk, reset => reset); --
    end block;
    -- CP-element group 607:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	605 
    -- CP-element group 607: successors 
    -- CP-element group 607: marked-successors 
    -- CP-element group 607: 	363 
    -- CP-element group 607: 	605 
    -- CP-element group 607:  members (3) 
      -- CP-element group 607: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/ra
      -- CP-element group 607: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/$exit
      -- CP-element group 607: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_sample_completed_
      -- 
    ra_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_0, ack => concat_CP_34_elements(607)); -- 
    -- CP-element group 608:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	606 
    -- CP-element group 608: successors 
    -- CP-element group 608: 	629 
    -- CP-element group 608: 	633 
    -- CP-element group 608: marked-successors 
    -- CP-element group 608: 	606 
    -- CP-element group 608:  members (3) 
      -- CP-element group 608: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/$exit
      -- CP-element group 608: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_update_completed_
      -- CP-element group 608: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/ca
      -- 
    ca_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 608_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_1, ack => concat_CP_34_elements(608)); -- 
    -- CP-element group 609:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	409 
    -- CP-element group 609: marked-predecessors 
    -- CP-element group 609: 	611 
    -- CP-element group 609: successors 
    -- CP-element group 609: 	611 
    -- CP-element group 609:  members (3) 
      -- CP-element group 609: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/$entry
      -- CP-element group 609: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/rr
      -- CP-element group 609: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_sample_start_
      -- 
    rr_2661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(609), ack => type_cast_1186_inst_req_0); -- 
    concat_cp_element_group_609: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_609"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(409) & concat_CP_34_elements(611);
      gj_concat_cp_element_group_609 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(609), clk => clk, reset => reset); --
    end block;
    -- CP-element group 610:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: marked-predecessors 
    -- CP-element group 610: 	612 
    -- CP-element group 610: 	615 
    -- CP-element group 610: 	675 
    -- CP-element group 610: successors 
    -- CP-element group 610: 	612 
    -- CP-element group 610:  members (3) 
      -- CP-element group 610: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_update_start_
      -- CP-element group 610: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/$entry
      -- CP-element group 610: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/cr
      -- 
    cr_2666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(610), ack => type_cast_1186_inst_req_1); -- 
    concat_cp_element_group_610: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_610"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(612) & concat_CP_34_elements(615) & concat_CP_34_elements(675);
      gj_concat_cp_element_group_610 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(610), clk => clk, reset => reset); --
    end block;
    -- CP-element group 611:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	609 
    -- CP-element group 611: successors 
    -- CP-element group 611: marked-successors 
    -- CP-element group 611: 	405 
    -- CP-element group 611: 	609 
    -- CP-element group 611:  members (3) 
      -- CP-element group 611: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/$exit
      -- CP-element group 611: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_sample_completed_
      -- CP-element group 611: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/ra
      -- 
    ra_2662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 611_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_0, ack => concat_CP_34_elements(611)); -- 
    -- CP-element group 612:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	610 
    -- CP-element group 612: successors 
    -- CP-element group 612: 	613 
    -- CP-element group 612: 	673 
    -- CP-element group 612: marked-successors 
    -- CP-element group 612: 	610 
    -- CP-element group 612:  members (3) 
      -- CP-element group 612: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_update_completed_
      -- CP-element group 612: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/$exit
      -- CP-element group 612: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/ca
      -- 
    ca_2667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 612_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_1, ack => concat_CP_34_elements(612)); -- 
    -- CP-element group 613:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	526 
    -- CP-element group 613: 	534 
    -- CP-element group 613: 	538 
    -- CP-element group 613: 	592 
    -- CP-element group 613: 	612 
    -- CP-element group 613: marked-predecessors 
    -- CP-element group 613: 	615 
    -- CP-element group 613: successors 
    -- CP-element group 613: 	615 
    -- CP-element group 613:  members (3) 
      -- CP-element group 613: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/$entry
      -- CP-element group 613: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/rr
      -- CP-element group 613: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_sample_start_
      -- 
    rr_2675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(613), ack => type_cast_1202_inst_req_0); -- 
    concat_cp_element_group_613: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_613"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(592) & concat_CP_34_elements(612) & concat_CP_34_elements(615);
      gj_concat_cp_element_group_613 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(613), clk => clk, reset => reset); --
    end block;
    -- CP-element group 614:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	319 
    -- CP-element group 614: marked-predecessors 
    -- CP-element group 614: 	616 
    -- CP-element group 614: 	687 
    -- CP-element group 614: successors 
    -- CP-element group 614: 	616 
    -- CP-element group 614:  members (3) 
      -- CP-element group 614: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_update_start_
      -- CP-element group 614: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/cr
      -- CP-element group 614: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/$entry
      -- 
    cr_2680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(614), ack => type_cast_1202_inst_req_1); -- 
    concat_cp_element_group_614: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_614"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(616) & concat_CP_34_elements(687);
      gj_concat_cp_element_group_614 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(614), clk => clk, reset => reset); --
    end block;
    -- CP-element group 615:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	613 
    -- CP-element group 615: successors 
    -- CP-element group 615: marked-successors 
    -- CP-element group 615: 	524 
    -- CP-element group 615: 	532 
    -- CP-element group 615: 	536 
    -- CP-element group 615: 	590 
    -- CP-element group 615: 	610 
    -- CP-element group 615: 	613 
    -- CP-element group 615:  members (3) 
      -- CP-element group 615: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/$exit
      -- CP-element group 615: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_sample_completed_
      -- CP-element group 615: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/ra
      -- 
    ra_2676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1202_inst_ack_0, ack => concat_CP_34_elements(615)); -- 
    -- CP-element group 616:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	614 
    -- CP-element group 616: successors 
    -- CP-element group 616: 	685 
    -- CP-element group 616: marked-successors 
    -- CP-element group 616: 	362 
    -- CP-element group 616: 	383 
    -- CP-element group 616: 	404 
    -- CP-element group 616: 	614 
    -- CP-element group 616: 	322 
    -- CP-element group 616:  members (3) 
      -- CP-element group 616: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_update_completed_
      -- CP-element group 616: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/ca
      -- CP-element group 616: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/$exit
      -- 
    ca_2681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 616_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1202_inst_ack_1, ack => concat_CP_34_elements(616)); -- 
    -- CP-element group 617:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	526 
    -- CP-element group 617: 	534 
    -- CP-element group 617: 	538 
    -- CP-element group 617: marked-predecessors 
    -- CP-element group 617: 	619 
    -- CP-element group 617: successors 
    -- CP-element group 617: 	619 
    -- CP-element group 617:  members (3) 
      -- CP-element group 617: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/req
      -- CP-element group 617: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/$entry
      -- CP-element group 617: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_sample_start_
      -- 
    req_2689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(617), ack => W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_req_0); -- 
    concat_cp_element_group_617: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_617"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(619);
      gj_concat_cp_element_group_617 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(617), clk => clk, reset => reset); --
    end block;
    -- CP-element group 618:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: marked-predecessors 
    -- CP-element group 618: 	620 
    -- CP-element group 618: successors 
    -- CP-element group 618: 	620 
    -- CP-element group 618:  members (3) 
      -- CP-element group 618: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/req
      -- CP-element group 618: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_update_start_
      -- 
    req_2694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(618), ack => W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_req_1); -- 
    concat_cp_element_group_618: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_618"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(620);
      gj_concat_cp_element_group_618 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(618), clk => clk, reset => reset); --
    end block;
    -- CP-element group 619:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	617 
    -- CP-element group 619: successors 
    -- CP-element group 619: marked-successors 
    -- CP-element group 619: 	524 
    -- CP-element group 619: 	532 
    -- CP-element group 619: 	536 
    -- CP-element group 619: 	617 
    -- CP-element group 619:  members (3) 
      -- CP-element group 619: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/ack
      -- CP-element group 619: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/$exit
      -- CP-element group 619: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_sample_completed_
      -- 
    ack_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 619_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_ack_0, ack => concat_CP_34_elements(619)); -- 
    -- CP-element group 620:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	618 
    -- CP-element group 620: successors 
    -- CP-element group 620: 	691 
    -- CP-element group 620: marked-successors 
    -- CP-element group 620: 	618 
    -- CP-element group 620:  members (3) 
      -- CP-element group 620: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/ack
      -- CP-element group 620: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_update_completed_
      -- CP-element group 620: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/$exit
      -- 
    ack_2695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 620_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_ack_1, ack => concat_CP_34_elements(620)); -- 
    -- CP-element group 621:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	526 
    -- CP-element group 621: 	534 
    -- CP-element group 621: 	538 
    -- CP-element group 621: marked-predecessors 
    -- CP-element group 621: 	623 
    -- CP-element group 621: successors 
    -- CP-element group 621: 	623 
    -- CP-element group 621:  members (3) 
      -- CP-element group 621: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_sample_start_
      -- CP-element group 621: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/$entry
      -- CP-element group 621: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/req
      -- 
    req_2703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(621), ack => W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_req_0); -- 
    concat_cp_element_group_621: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_621"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(623);
      gj_concat_cp_element_group_621 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(621), clk => clk, reset => reset); --
    end block;
    -- CP-element group 622:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	319 
    -- CP-element group 622: marked-predecessors 
    -- CP-element group 622: 	624 
    -- CP-element group 622: 	687 
    -- CP-element group 622: successors 
    -- CP-element group 622: 	624 
    -- CP-element group 622:  members (3) 
      -- CP-element group 622: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/req
      -- CP-element group 622: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_update_start_
      -- CP-element group 622: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/$entry
      -- 
    req_2708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(622), ack => W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_req_1); -- 
    concat_cp_element_group_622: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_622"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(624) & concat_CP_34_elements(687);
      gj_concat_cp_element_group_622 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(622), clk => clk, reset => reset); --
    end block;
    -- CP-element group 623:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	621 
    -- CP-element group 623: successors 
    -- CP-element group 623: marked-successors 
    -- CP-element group 623: 	524 
    -- CP-element group 623: 	532 
    -- CP-element group 623: 	536 
    -- CP-element group 623: 	621 
    -- CP-element group 623:  members (3) 
      -- CP-element group 623: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_sample_completed_
      -- CP-element group 623: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/$exit
      -- CP-element group 623: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/ack
      -- 
    ack_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 623_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_ack_0, ack => concat_CP_34_elements(623)); -- 
    -- CP-element group 624:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	622 
    -- CP-element group 624: successors 
    -- CP-element group 624: 	685 
    -- CP-element group 624: marked-successors 
    -- CP-element group 624: 	362 
    -- CP-element group 624: 	383 
    -- CP-element group 624: 	404 
    -- CP-element group 624: 	622 
    -- CP-element group 624: 	322 
    -- CP-element group 624:  members (3) 
      -- CP-element group 624: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/$exit
      -- CP-element group 624: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/ack
      -- CP-element group 624: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_update_completed_
      -- 
    ack_2709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 624_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_ack_1, ack => concat_CP_34_elements(624)); -- 
    -- CP-element group 625:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	526 
    -- CP-element group 625: 	534 
    -- CP-element group 625: 	538 
    -- CP-element group 625: marked-predecessors 
    -- CP-element group 625: 	627 
    -- CP-element group 625: successors 
    -- CP-element group 625: 	627 
    -- CP-element group 625:  members (3) 
      -- CP-element group 625: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/req
      -- CP-element group 625: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/$entry
      -- CP-element group 625: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_sample_start_
      -- 
    req_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(625), ack => W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_req_0); -- 
    concat_cp_element_group_625: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_625"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(627);
      gj_concat_cp_element_group_625 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(625), clk => clk, reset => reset); --
    end block;
    -- CP-element group 626:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	319 
    -- CP-element group 626: marked-predecessors 
    -- CP-element group 626: 	628 
    -- CP-element group 626: 	687 
    -- CP-element group 626: successors 
    -- CP-element group 626: 	628 
    -- CP-element group 626:  members (3) 
      -- CP-element group 626: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/req
      -- CP-element group 626: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/$entry
      -- CP-element group 626: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_update_start_
      -- 
    req_2722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(626), ack => W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_req_1); -- 
    concat_cp_element_group_626: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_626"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(628) & concat_CP_34_elements(687);
      gj_concat_cp_element_group_626 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(626), clk => clk, reset => reset); --
    end block;
    -- CP-element group 627:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	625 
    -- CP-element group 627: successors 
    -- CP-element group 627: marked-successors 
    -- CP-element group 627: 	524 
    -- CP-element group 627: 	532 
    -- CP-element group 627: 	536 
    -- CP-element group 627: 	625 
    -- CP-element group 627:  members (3) 
      -- CP-element group 627: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/ack
      -- CP-element group 627: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/$exit
      -- CP-element group 627: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_sample_completed_
      -- 
    ack_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_ack_0, ack => concat_CP_34_elements(627)); -- 
    -- CP-element group 628:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	626 
    -- CP-element group 628: successors 
    -- CP-element group 628: 	685 
    -- CP-element group 628: marked-successors 
    -- CP-element group 628: 	362 
    -- CP-element group 628: 	383 
    -- CP-element group 628: 	404 
    -- CP-element group 628: 	626 
    -- CP-element group 628: 	322 
    -- CP-element group 628:  members (3) 
      -- CP-element group 628: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/ack
      -- CP-element group 628: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/$exit
      -- CP-element group 628: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_update_completed_
      -- 
    ack_2723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 628_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_ack_1, ack => concat_CP_34_elements(628)); -- 
    -- CP-element group 629:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	526 
    -- CP-element group 629: 	534 
    -- CP-element group 629: 	538 
    -- CP-element group 629: 	596 
    -- CP-element group 629: 	608 
    -- CP-element group 629: marked-predecessors 
    -- CP-element group 629: 	631 
    -- CP-element group 629: successors 
    -- CP-element group 629: 	631 
    -- CP-element group 629:  members (3) 
      -- CP-element group 629: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/rr
      -- CP-element group 629: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_sample_start_
      -- CP-element group 629: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/$entry
      -- 
    rr_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(629), ack => type_cast_1238_inst_req_0); -- 
    concat_cp_element_group_629: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_629"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(596) & concat_CP_34_elements(608) & concat_CP_34_elements(631);
      gj_concat_cp_element_group_629 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(629), clk => clk, reset => reset); --
    end block;
    -- CP-element group 630:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	319 
    -- CP-element group 630: marked-predecessors 
    -- CP-element group 630: 	632 
    -- CP-element group 630: successors 
    -- CP-element group 630: 	632 
    -- CP-element group 630:  members (3) 
      -- CP-element group 630: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_update_start_
      -- CP-element group 630: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/$entry
      -- CP-element group 630: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/cr
      -- 
    cr_2736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(630), ack => type_cast_1238_inst_req_1); -- 
    concat_cp_element_group_630: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_630"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(632);
      gj_concat_cp_element_group_630 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(630), clk => clk, reset => reset); --
    end block;
    -- CP-element group 631:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	629 
    -- CP-element group 631: successors 
    -- CP-element group 631: marked-successors 
    -- CP-element group 631: 	524 
    -- CP-element group 631: 	532 
    -- CP-element group 631: 	536 
    -- CP-element group 631: 	594 
    -- CP-element group 631: 	606 
    -- CP-element group 631: 	629 
    -- CP-element group 631:  members (3) 
      -- CP-element group 631: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/ra
      -- CP-element group 631: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_sample_completed_
      -- CP-element group 631: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/$exit
      -- 
    ra_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 631_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => concat_CP_34_elements(631)); -- 
    -- CP-element group 632:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	630 
    -- CP-element group 632: successors 
    -- CP-element group 632: 	691 
    -- CP-element group 632: marked-successors 
    -- CP-element group 632: 	362 
    -- CP-element group 632: 	630 
    -- CP-element group 632:  members (3) 
      -- CP-element group 632: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_update_completed_
      -- CP-element group 632: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/$exit
      -- CP-element group 632: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/ca
      -- 
    ca_2737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 632_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => concat_CP_34_elements(632)); -- 
    -- CP-element group 633:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	526 
    -- CP-element group 633: 	534 
    -- CP-element group 633: 	538 
    -- CP-element group 633: 	596 
    -- CP-element group 633: 	608 
    -- CP-element group 633: marked-predecessors 
    -- CP-element group 633: 	635 
    -- CP-element group 633: successors 
    -- CP-element group 633: 	635 
    -- CP-element group 633:  members (3) 
      -- CP-element group 633: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_sample_start_
      -- CP-element group 633: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/$entry
      -- CP-element group 633: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/rr
      -- 
    rr_2745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(633), ack => type_cast_1242_inst_req_0); -- 
    concat_cp_element_group_633: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_633"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(596) & concat_CP_34_elements(608) & concat_CP_34_elements(635);
      gj_concat_cp_element_group_633 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(633), clk => clk, reset => reset); --
    end block;
    -- CP-element group 634:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	319 
    -- CP-element group 634: marked-predecessors 
    -- CP-element group 634: 	636 
    -- CP-element group 634: successors 
    -- CP-element group 634: 	636 
    -- CP-element group 634:  members (3) 
      -- CP-element group 634: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_update_start_
      -- CP-element group 634: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/$entry
      -- CP-element group 634: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/cr
      -- 
    cr_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(634), ack => type_cast_1242_inst_req_1); -- 
    concat_cp_element_group_634: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_634"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(636);
      gj_concat_cp_element_group_634 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(634), clk => clk, reset => reset); --
    end block;
    -- CP-element group 635:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	633 
    -- CP-element group 635: successors 
    -- CP-element group 635: marked-successors 
    -- CP-element group 635: 	524 
    -- CP-element group 635: 	532 
    -- CP-element group 635: 	536 
    -- CP-element group 635: 	594 
    -- CP-element group 635: 	606 
    -- CP-element group 635: 	633 
    -- CP-element group 635:  members (3) 
      -- CP-element group 635: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/$exit
      -- CP-element group 635: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_sample_completed_
      -- CP-element group 635: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/ra
      -- 
    ra_2746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_0, ack => concat_CP_34_elements(635)); -- 
    -- CP-element group 636:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	634 
    -- CP-element group 636: successors 
    -- CP-element group 636: 	691 
    -- CP-element group 636: marked-successors 
    -- CP-element group 636: 	362 
    -- CP-element group 636: 	634 
    -- CP-element group 636:  members (3) 
      -- CP-element group 636: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_update_completed_
      -- CP-element group 636: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/$exit
      -- CP-element group 636: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/ca
      -- 
    ca_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 636_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_1, ack => concat_CP_34_elements(636)); -- 
    -- CP-element group 637:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	367 
    -- CP-element group 637: marked-predecessors 
    -- CP-element group 637: 	639 
    -- CP-element group 637: successors 
    -- CP-element group 637: 	639 
    -- CP-element group 637:  members (3) 
      -- CP-element group 637: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_sample_start_
      -- CP-element group 637: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/$entry
      -- CP-element group 637: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/rr
      -- 
    rr_2759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(637), ack => type_cast_1246_inst_req_0); -- 
    concat_cp_element_group_637: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_637"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(367) & concat_CP_34_elements(639);
      gj_concat_cp_element_group_637 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(637), clk => clk, reset => reset); --
    end block;
    -- CP-element group 638:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: marked-predecessors 
    -- CP-element group 638: 	640 
    -- CP-element group 638: 	643 
    -- CP-element group 638: successors 
    -- CP-element group 638: 	640 
    -- CP-element group 638:  members (3) 
      -- CP-element group 638: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_update_start_
      -- CP-element group 638: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/cr
      -- 
    cr_2764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(638), ack => type_cast_1246_inst_req_1); -- 
    concat_cp_element_group_638: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_638"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(640) & concat_CP_34_elements(643);
      gj_concat_cp_element_group_638 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(638), clk => clk, reset => reset); --
    end block;
    -- CP-element group 639:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	637 
    -- CP-element group 639: successors 
    -- CP-element group 639: marked-successors 
    -- CP-element group 639: 	363 
    -- CP-element group 639: 	637 
    -- CP-element group 639:  members (3) 
      -- CP-element group 639: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_sample_completed_
      -- CP-element group 639: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/$exit
      -- CP-element group 639: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/ra
      -- 
    ra_2760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 639_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_0, ack => concat_CP_34_elements(639)); -- 
    -- CP-element group 640:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	638 
    -- CP-element group 640: successors 
    -- CP-element group 640: 	641 
    -- CP-element group 640: marked-successors 
    -- CP-element group 640: 	638 
    -- CP-element group 640:  members (3) 
      -- CP-element group 640: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_update_completed_
      -- CP-element group 640: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/$exit
      -- CP-element group 640: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/ca
      -- 
    ca_2765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 640_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_1, ack => concat_CP_34_elements(640)); -- 
    -- CP-element group 641:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	506 
    -- CP-element group 641: 	518 
    -- CP-element group 641: 	640 
    -- CP-element group 641: marked-predecessors 
    -- CP-element group 641: 	643 
    -- CP-element group 641: successors 
    -- CP-element group 641: 	643 
    -- CP-element group 641:  members (3) 
      -- CP-element group 641: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/req
      -- CP-element group 641: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_sample_start_
      -- CP-element group 641: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/$entry
      -- 
    req_2773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(641), ack => MUX_1253_inst_req_0); -- 
    concat_cp_element_group_641: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_641"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(518) & concat_CP_34_elements(640) & concat_CP_34_elements(643);
      gj_concat_cp_element_group_641 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(641), clk => clk, reset => reset); --
    end block;
    -- CP-element group 642:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	319 
    -- CP-element group 642: marked-predecessors 
    -- CP-element group 642: 	644 
    -- CP-element group 642: successors 
    -- CP-element group 642: 	644 
    -- CP-element group 642:  members (3) 
      -- CP-element group 642: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/$entry
      -- CP-element group 642: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_update_start_
      -- CP-element group 642: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/req
      -- 
    req_2778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(642), ack => MUX_1253_inst_req_1); -- 
    concat_cp_element_group_642: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_642"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(644);
      gj_concat_cp_element_group_642 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(642), clk => clk, reset => reset); --
    end block;
    -- CP-element group 643:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	641 
    -- CP-element group 643: successors 
    -- CP-element group 643: marked-successors 
    -- CP-element group 643: 	504 
    -- CP-element group 643: 	516 
    -- CP-element group 643: 	638 
    -- CP-element group 643: 	641 
    -- CP-element group 643:  members (3) 
      -- CP-element group 643: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_sample_completed_
      -- CP-element group 643: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/$exit
      -- CP-element group 643: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/ack
      -- 
    ack_2774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 643_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1253_inst_ack_0, ack => concat_CP_34_elements(643)); -- 
    -- CP-element group 644:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	642 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	691 
    -- CP-element group 644: marked-successors 
    -- CP-element group 644: 	362 
    -- CP-element group 644: 	642 
    -- CP-element group 644:  members (3) 
      -- CP-element group 644: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/ack
      -- CP-element group 644: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/$exit
      -- CP-element group 644: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_update_completed_
      -- 
    ack_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 644_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1253_inst_ack_1, ack => concat_CP_34_elements(644)); -- 
    -- CP-element group 645:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	526 
    -- CP-element group 645: 	534 
    -- CP-element group 645: 	538 
    -- CP-element group 645: 	600 
    -- CP-element group 645: 	604 
    -- CP-element group 645: marked-predecessors 
    -- CP-element group 645: 	647 
    -- CP-element group 645: successors 
    -- CP-element group 645: 	647 
    -- CP-element group 645:  members (3) 
      -- CP-element group 645: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_sample_start_
      -- CP-element group 645: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/$entry
      -- CP-element group 645: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/rr
      -- 
    rr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(645), ack => type_cast_1266_inst_req_0); -- 
    concat_cp_element_group_645: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_645"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(600) & concat_CP_34_elements(604) & concat_CP_34_elements(647);
      gj_concat_cp_element_group_645 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(645), clk => clk, reset => reset); --
    end block;
    -- CP-element group 646:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	319 
    -- CP-element group 646: marked-predecessors 
    -- CP-element group 646: 	648 
    -- CP-element group 646: 	687 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	648 
    -- CP-element group 646:  members (3) 
      -- CP-element group 646: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_update_start_
      -- CP-element group 646: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/$entry
      -- CP-element group 646: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/cr
      -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(646), ack => type_cast_1266_inst_req_1); -- 
    concat_cp_element_group_646: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_646"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(648) & concat_CP_34_elements(687);
      gj_concat_cp_element_group_646 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(646), clk => clk, reset => reset); --
    end block;
    -- CP-element group 647:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	645 
    -- CP-element group 647: successors 
    -- CP-element group 647: marked-successors 
    -- CP-element group 647: 	524 
    -- CP-element group 647: 	532 
    -- CP-element group 647: 	536 
    -- CP-element group 647: 	598 
    -- CP-element group 647: 	602 
    -- CP-element group 647: 	645 
    -- CP-element group 647:  members (3) 
      -- CP-element group 647: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_sample_completed_
      -- CP-element group 647: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/$exit
      -- CP-element group 647: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/ra
      -- 
    ra_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 647_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_0, ack => concat_CP_34_elements(647)); -- 
    -- CP-element group 648:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	646 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	685 
    -- CP-element group 648: marked-successors 
    -- CP-element group 648: 	646 
    -- CP-element group 648: 	322 
    -- CP-element group 648:  members (3) 
      -- CP-element group 648: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_update_completed_
      -- CP-element group 648: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/$exit
      -- CP-element group 648: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/ca
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 648_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_1, ack => concat_CP_34_elements(648)); -- 
    -- CP-element group 649:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	526 
    -- CP-element group 649: 	534 
    -- CP-element group 649: 	538 
    -- CP-element group 649: 	600 
    -- CP-element group 649: 	604 
    -- CP-element group 649: marked-predecessors 
    -- CP-element group 649: 	651 
    -- CP-element group 649: successors 
    -- CP-element group 649: 	651 
    -- CP-element group 649:  members (3) 
      -- CP-element group 649: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/rr
      -- CP-element group 649: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/$entry
      -- CP-element group 649: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_sample_start_
      -- 
    rr_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(649), ack => type_cast_1270_inst_req_0); -- 
    concat_cp_element_group_649: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_649"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(600) & concat_CP_34_elements(604) & concat_CP_34_elements(651);
      gj_concat_cp_element_group_649 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(649), clk => clk, reset => reset); --
    end block;
    -- CP-element group 650:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	319 
    -- CP-element group 650: marked-predecessors 
    -- CP-element group 650: 	652 
    -- CP-element group 650: 	687 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	652 
    -- CP-element group 650:  members (3) 
      -- CP-element group 650: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/$entry
      -- CP-element group 650: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/cr
      -- CP-element group 650: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_update_start_
      -- 
    cr_2806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(650), ack => type_cast_1270_inst_req_1); -- 
    concat_cp_element_group_650: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_650"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(652) & concat_CP_34_elements(687);
      gj_concat_cp_element_group_650 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(650), clk => clk, reset => reset); --
    end block;
    -- CP-element group 651:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	649 
    -- CP-element group 651: successors 
    -- CP-element group 651: marked-successors 
    -- CP-element group 651: 	524 
    -- CP-element group 651: 	532 
    -- CP-element group 651: 	536 
    -- CP-element group 651: 	598 
    -- CP-element group 651: 	602 
    -- CP-element group 651: 	649 
    -- CP-element group 651:  members (3) 
      -- CP-element group 651: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/$exit
      -- CP-element group 651: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/ra
      -- CP-element group 651: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_sample_completed_
      -- 
    ra_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 651_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_0, ack => concat_CP_34_elements(651)); -- 
    -- CP-element group 652:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	650 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	685 
    -- CP-element group 652: marked-successors 
    -- CP-element group 652: 	650 
    -- CP-element group 652: 	322 
    -- CP-element group 652:  members (3) 
      -- CP-element group 652: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_update_completed_
      -- CP-element group 652: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/ca
      -- CP-element group 652: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/$exit
      -- 
    ca_2807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 652_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_1, ack => concat_CP_34_elements(652)); -- 
    -- CP-element group 653:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	428 
    -- CP-element group 653: 	490 
    -- CP-element group 653: 	494 
    -- CP-element group 653: marked-predecessors 
    -- CP-element group 653: 	655 
    -- CP-element group 653: successors 
    -- CP-element group 653: 	655 
    -- CP-element group 653:  members (3) 
      -- CP-element group 653: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/$entry
      -- CP-element group 653: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/rr
      -- CP-element group 653: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_sample_start_
      -- 
    rr_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(653), ack => type_cast_1274_inst_req_0); -- 
    concat_cp_element_group_653: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_653"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(490) & concat_CP_34_elements(494) & concat_CP_34_elements(655);
      gj_concat_cp_element_group_653 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(653), clk => clk, reset => reset); --
    end block;
    -- CP-element group 654:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: marked-predecessors 
    -- CP-element group 654: 	656 
    -- CP-element group 654: 	659 
    -- CP-element group 654: successors 
    -- CP-element group 654: 	656 
    -- CP-element group 654:  members (3) 
      -- CP-element group 654: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_update_start_
      -- CP-element group 654: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/cr
      -- CP-element group 654: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/$entry
      -- 
    cr_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(654), ack => type_cast_1274_inst_req_1); -- 
    concat_cp_element_group_654: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_654"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(656) & concat_CP_34_elements(659);
      gj_concat_cp_element_group_654 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(654), clk => clk, reset => reset); --
    end block;
    -- CP-element group 655:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	653 
    -- CP-element group 655: successors 
    -- CP-element group 655: marked-successors 
    -- CP-element group 655: 	426 
    -- CP-element group 655: 	488 
    -- CP-element group 655: 	492 
    -- CP-element group 655: 	653 
    -- CP-element group 655:  members (3) 
      -- CP-element group 655: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/ra
      -- CP-element group 655: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_sample_completed_
      -- CP-element group 655: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/$exit
      -- 
    ra_2816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 655_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_0, ack => concat_CP_34_elements(655)); -- 
    -- CP-element group 656:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	654 
    -- CP-element group 656: successors 
    -- CP-element group 656: 	657 
    -- CP-element group 656: marked-successors 
    -- CP-element group 656: 	654 
    -- CP-element group 656:  members (3) 
      -- CP-element group 656: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_update_completed_
      -- CP-element group 656: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/$exit
      -- CP-element group 656: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/ca
      -- 
    ca_2821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 656_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_1, ack => concat_CP_34_elements(656)); -- 
    -- CP-element group 657:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	506 
    -- CP-element group 657: 	518 
    -- CP-element group 657: 	656 
    -- CP-element group 657: marked-predecessors 
    -- CP-element group 657: 	659 
    -- CP-element group 657: successors 
    -- CP-element group 657: 	659 
    -- CP-element group 657:  members (3) 
      -- CP-element group 657: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_sample_start_
      -- CP-element group 657: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/$entry
      -- CP-element group 657: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/req
      -- 
    req_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(657), ack => MUX_1281_inst_req_0); -- 
    concat_cp_element_group_657: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_657"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(518) & concat_CP_34_elements(656) & concat_CP_34_elements(659);
      gj_concat_cp_element_group_657 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(657), clk => clk, reset => reset); --
    end block;
    -- CP-element group 658:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	319 
    -- CP-element group 658: marked-predecessors 
    -- CP-element group 658: 	660 
    -- CP-element group 658: 	687 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	660 
    -- CP-element group 658:  members (3) 
      -- CP-element group 658: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_update_start_
      -- CP-element group 658: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/$entry
      -- CP-element group 658: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/req
      -- 
    req_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(658), ack => MUX_1281_inst_req_1); -- 
    concat_cp_element_group_658: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_658"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(660) & concat_CP_34_elements(687);
      gj_concat_cp_element_group_658 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(658), clk => clk, reset => reset); --
    end block;
    -- CP-element group 659:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	657 
    -- CP-element group 659: successors 
    -- CP-element group 659: marked-successors 
    -- CP-element group 659: 	504 
    -- CP-element group 659: 	516 
    -- CP-element group 659: 	654 
    -- CP-element group 659: 	657 
    -- CP-element group 659:  members (3) 
      -- CP-element group 659: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_sample_completed_
      -- CP-element group 659: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/$exit
      -- CP-element group 659: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/ack
      -- 
    ack_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 659_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1281_inst_ack_0, ack => concat_CP_34_elements(659)); -- 
    -- CP-element group 660:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	658 
    -- CP-element group 660: successors 
    -- CP-element group 660: 	685 
    -- CP-element group 660: marked-successors 
    -- CP-element group 660: 	658 
    -- CP-element group 660: 	322 
    -- CP-element group 660:  members (3) 
      -- CP-element group 660: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_update_completed_
      -- CP-element group 660: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/$exit
      -- CP-element group 660: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/ack
      -- 
    ack_2835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 660_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1281_inst_ack_1, ack => concat_CP_34_elements(660)); -- 
    -- CP-element group 661:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	428 
    -- CP-element group 661: 	482 
    -- CP-element group 661: 	502 
    -- CP-element group 661: marked-predecessors 
    -- CP-element group 661: 	663 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	663 
    -- CP-element group 661:  members (3) 
      -- CP-element group 661: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_sample_start_
      -- CP-element group 661: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/$entry
      -- CP-element group 661: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/rr
      -- 
    rr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(661), ack => type_cast_1294_inst_req_0); -- 
    concat_cp_element_group_661: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_661"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(482) & concat_CP_34_elements(502) & concat_CP_34_elements(663);
      gj_concat_cp_element_group_661 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(661), clk => clk, reset => reset); --
    end block;
    -- CP-element group 662:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	319 
    -- CP-element group 662: marked-predecessors 
    -- CP-element group 662: 	664 
    -- CP-element group 662: successors 
    -- CP-element group 662: 	664 
    -- CP-element group 662:  members (3) 
      -- CP-element group 662: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_update_start_
      -- CP-element group 662: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/$entry
      -- CP-element group 662: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/cr
      -- 
    cr_2848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(662), ack => type_cast_1294_inst_req_1); -- 
    concat_cp_element_group_662: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_662"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(664);
      gj_concat_cp_element_group_662 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(662), clk => clk, reset => reset); --
    end block;
    -- CP-element group 663:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	661 
    -- CP-element group 663: successors 
    -- CP-element group 663: marked-successors 
    -- CP-element group 663: 	426 
    -- CP-element group 663: 	480 
    -- CP-element group 663: 	500 
    -- CP-element group 663: 	661 
    -- CP-element group 663:  members (3) 
      -- CP-element group 663: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_sample_completed_
      -- CP-element group 663: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/$exit
      -- CP-element group 663: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/ra
      -- 
    ra_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1294_inst_ack_0, ack => concat_CP_34_elements(663)); -- 
    -- CP-element group 664:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	662 
    -- CP-element group 664: successors 
    -- CP-element group 664: 	691 
    -- CP-element group 664: marked-successors 
    -- CP-element group 664: 	383 
    -- CP-element group 664: 	662 
    -- CP-element group 664:  members (3) 
      -- CP-element group 664: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_update_completed_
      -- CP-element group 664: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/$exit
      -- CP-element group 664: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/ca
      -- 
    ca_2849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 664_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1294_inst_ack_1, ack => concat_CP_34_elements(664)); -- 
    -- CP-element group 665:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	428 
    -- CP-element group 665: 	482 
    -- CP-element group 665: 	502 
    -- CP-element group 665: marked-predecessors 
    -- CP-element group 665: 	667 
    -- CP-element group 665: successors 
    -- CP-element group 665: 	667 
    -- CP-element group 665:  members (3) 
      -- CP-element group 665: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_sample_start_
      -- CP-element group 665: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/$entry
      -- CP-element group 665: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/rr
      -- 
    rr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(665), ack => type_cast_1298_inst_req_0); -- 
    concat_cp_element_group_665: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_665"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(428) & concat_CP_34_elements(482) & concat_CP_34_elements(502) & concat_CP_34_elements(667);
      gj_concat_cp_element_group_665 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(665), clk => clk, reset => reset); --
    end block;
    -- CP-element group 666:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: marked-predecessors 
    -- CP-element group 666: 	668 
    -- CP-element group 666: 	671 
    -- CP-element group 666: successors 
    -- CP-element group 666: 	668 
    -- CP-element group 666:  members (3) 
      -- CP-element group 666: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/cr
      -- 
    cr_2862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_1298_inst_req_1); -- 
    concat_cp_element_group_666: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_666"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(668) & concat_CP_34_elements(671);
      gj_concat_cp_element_group_666 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(666), clk => clk, reset => reset); --
    end block;
    -- CP-element group 667:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	665 
    -- CP-element group 667: successors 
    -- CP-element group 667: marked-successors 
    -- CP-element group 667: 	426 
    -- CP-element group 667: 	480 
    -- CP-element group 667: 	500 
    -- CP-element group 667: 	665 
    -- CP-element group 667:  members (3) 
      -- CP-element group 667: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_sample_completed_
      -- CP-element group 667: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/$exit
      -- CP-element group 667: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/ra
      -- 
    ra_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 667_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1298_inst_ack_0, ack => concat_CP_34_elements(667)); -- 
    -- CP-element group 668:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	666 
    -- CP-element group 668: successors 
    -- CP-element group 668: 	669 
    -- CP-element group 668: marked-successors 
    -- CP-element group 668: 	666 
    -- CP-element group 668:  members (3) 
      -- CP-element group 668: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_update_completed_
      -- CP-element group 668: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/$exit
      -- CP-element group 668: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/ca
      -- 
    ca_2863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 668_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1298_inst_ack_1, ack => concat_CP_34_elements(668)); -- 
    -- CP-element group 669:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	506 
    -- CP-element group 669: 	518 
    -- CP-element group 669: 	668 
    -- CP-element group 669: marked-predecessors 
    -- CP-element group 669: 	671 
    -- CP-element group 669: successors 
    -- CP-element group 669: 	671 
    -- CP-element group 669:  members (3) 
      -- CP-element group 669: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_sample_start_
      -- CP-element group 669: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/$entry
      -- CP-element group 669: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/req
      -- 
    req_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(669), ack => MUX_1305_inst_req_0); -- 
    concat_cp_element_group_669: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_669"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(518) & concat_CP_34_elements(668) & concat_CP_34_elements(671);
      gj_concat_cp_element_group_669 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(669), clk => clk, reset => reset); --
    end block;
    -- CP-element group 670:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	319 
    -- CP-element group 670: marked-predecessors 
    -- CP-element group 670: 	672 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	672 
    -- CP-element group 670:  members (3) 
      -- CP-element group 670: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_update_start_
      -- CP-element group 670: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/$entry
      -- CP-element group 670: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/req
      -- 
    req_2876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(670), ack => MUX_1305_inst_req_1); -- 
    concat_cp_element_group_670: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_670"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(672);
      gj_concat_cp_element_group_670 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(670), clk => clk, reset => reset); --
    end block;
    -- CP-element group 671:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	669 
    -- CP-element group 671: successors 
    -- CP-element group 671: marked-successors 
    -- CP-element group 671: 	504 
    -- CP-element group 671: 	516 
    -- CP-element group 671: 	666 
    -- CP-element group 671: 	669 
    -- CP-element group 671:  members (3) 
      -- CP-element group 671: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_sample_completed_
      -- CP-element group 671: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/$exit
      -- CP-element group 671: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/ack
      -- 
    ack_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 671_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1305_inst_ack_0, ack => concat_CP_34_elements(671)); -- 
    -- CP-element group 672:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	670 
    -- CP-element group 672: successors 
    -- CP-element group 672: 	691 
    -- CP-element group 672: marked-successors 
    -- CP-element group 672: 	383 
    -- CP-element group 672: 	670 
    -- CP-element group 672:  members (3) 
      -- CP-element group 672: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_update_completed_
      -- CP-element group 672: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/$exit
      -- CP-element group 672: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/ack
      -- 
    ack_2877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 672_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1305_inst_ack_1, ack => concat_CP_34_elements(672)); -- 
    -- CP-element group 673:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	526 
    -- CP-element group 673: 	534 
    -- CP-element group 673: 	538 
    -- CP-element group 673: 	592 
    -- CP-element group 673: 	612 
    -- CP-element group 673: marked-predecessors 
    -- CP-element group 673: 	675 
    -- CP-element group 673: successors 
    -- CP-element group 673: 	675 
    -- CP-element group 673:  members (3) 
      -- CP-element group 673: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_sample_start_
      -- CP-element group 673: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/rr
      -- 
    rr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1320_inst_req_0); -- 
    concat_cp_element_group_673: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_673"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(526) & concat_CP_34_elements(534) & concat_CP_34_elements(538) & concat_CP_34_elements(592) & concat_CP_34_elements(612) & concat_CP_34_elements(675);
      gj_concat_cp_element_group_673 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(673), clk => clk, reset => reset); --
    end block;
    -- CP-element group 674:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	319 
    -- CP-element group 674: marked-predecessors 
    -- CP-element group 674: 	676 
    -- CP-element group 674: successors 
    -- CP-element group 674: 	676 
    -- CP-element group 674:  members (3) 
      -- CP-element group 674: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_update_start_
      -- CP-element group 674: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/$entry
      -- CP-element group 674: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/cr
      -- 
    cr_2890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(674), ack => type_cast_1320_inst_req_1); -- 
    concat_cp_element_group_674: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_674"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(676);
      gj_concat_cp_element_group_674 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(674), clk => clk, reset => reset); --
    end block;
    -- CP-element group 675:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 675: predecessors 
    -- CP-element group 675: 	673 
    -- CP-element group 675: successors 
    -- CP-element group 675: marked-successors 
    -- CP-element group 675: 	524 
    -- CP-element group 675: 	532 
    -- CP-element group 675: 	536 
    -- CP-element group 675: 	590 
    -- CP-element group 675: 	610 
    -- CP-element group 675: 	673 
    -- CP-element group 675:  members (3) 
      -- CP-element group 675: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_sample_completed_
      -- CP-element group 675: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/$exit
      -- CP-element group 675: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/ra
      -- 
    ra_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 675_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_0, ack => concat_CP_34_elements(675)); -- 
    -- CP-element group 676:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 676: predecessors 
    -- CP-element group 676: 	674 
    -- CP-element group 676: successors 
    -- CP-element group 676: 	691 
    -- CP-element group 676: marked-successors 
    -- CP-element group 676: 	404 
    -- CP-element group 676: 	674 
    -- CP-element group 676:  members (3) 
      -- CP-element group 676: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_update_completed_
      -- CP-element group 676: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/$exit
      -- CP-element group 676: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/ca
      -- 
    ca_2891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 676_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_1, ack => concat_CP_34_elements(676)); -- 
    -- CP-element group 677:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 677: predecessors 
    -- CP-element group 677: 	409 
    -- CP-element group 677: marked-predecessors 
    -- CP-element group 677: 	679 
    -- CP-element group 677: successors 
    -- CP-element group 677: 	679 
    -- CP-element group 677:  members (3) 
      -- CP-element group 677: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_sample_start_
      -- CP-element group 677: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/$entry
      -- CP-element group 677: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/rr
      -- 
    rr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(677), ack => type_cast_1324_inst_req_0); -- 
    concat_cp_element_group_677: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_677"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(409) & concat_CP_34_elements(679);
      gj_concat_cp_element_group_677 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(677), clk => clk, reset => reset); --
    end block;
    -- CP-element group 678:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 678: predecessors 
    -- CP-element group 678: marked-predecessors 
    -- CP-element group 678: 	680 
    -- CP-element group 678: 	683 
    -- CP-element group 678: successors 
    -- CP-element group 678: 	680 
    -- CP-element group 678:  members (3) 
      -- CP-element group 678: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_update_start_
      -- CP-element group 678: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/$entry
      -- CP-element group 678: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/cr
      -- 
    cr_2904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(678), ack => type_cast_1324_inst_req_1); -- 
    concat_cp_element_group_678: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_678"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(680) & concat_CP_34_elements(683);
      gj_concat_cp_element_group_678 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(678), clk => clk, reset => reset); --
    end block;
    -- CP-element group 679:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 679: predecessors 
    -- CP-element group 679: 	677 
    -- CP-element group 679: successors 
    -- CP-element group 679: marked-successors 
    -- CP-element group 679: 	405 
    -- CP-element group 679: 	677 
    -- CP-element group 679:  members (3) 
      -- CP-element group 679: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_sample_completed_
      -- CP-element group 679: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/$exit
      -- CP-element group 679: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/ra
      -- 
    ra_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 679_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1324_inst_ack_0, ack => concat_CP_34_elements(679)); -- 
    -- CP-element group 680:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 680: predecessors 
    -- CP-element group 680: 	678 
    -- CP-element group 680: successors 
    -- CP-element group 680: 	681 
    -- CP-element group 680: marked-successors 
    -- CP-element group 680: 	678 
    -- CP-element group 680:  members (3) 
      -- CP-element group 680: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_update_completed_
      -- CP-element group 680: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/$exit
      -- CP-element group 680: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/ca
      -- 
    ca_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 680_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1324_inst_ack_1, ack => concat_CP_34_elements(680)); -- 
    -- CP-element group 681:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 681: predecessors 
    -- CP-element group 681: 	506 
    -- CP-element group 681: 	518 
    -- CP-element group 681: 	680 
    -- CP-element group 681: marked-predecessors 
    -- CP-element group 681: 	683 
    -- CP-element group 681: successors 
    -- CP-element group 681: 	683 
    -- CP-element group 681:  members (3) 
      -- CP-element group 681: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_sample_start_
      -- CP-element group 681: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/$entry
      -- CP-element group 681: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/req
      -- 
    req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(681), ack => MUX_1331_inst_req_0); -- 
    concat_cp_element_group_681: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_681"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(506) & concat_CP_34_elements(518) & concat_CP_34_elements(680) & concat_CP_34_elements(683);
      gj_concat_cp_element_group_681 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(681), clk => clk, reset => reset); --
    end block;
    -- CP-element group 682:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 682: predecessors 
    -- CP-element group 682: 	319 
    -- CP-element group 682: marked-predecessors 
    -- CP-element group 682: 	684 
    -- CP-element group 682: successors 
    -- CP-element group 682: 	684 
    -- CP-element group 682:  members (3) 
      -- CP-element group 682: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_update_start_
      -- CP-element group 682: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/$entry
      -- CP-element group 682: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/req
      -- 
    req_2918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(682), ack => MUX_1331_inst_req_1); -- 
    concat_cp_element_group_682: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_682"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(684);
      gj_concat_cp_element_group_682 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(682), clk => clk, reset => reset); --
    end block;
    -- CP-element group 683:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 683: predecessors 
    -- CP-element group 683: 	681 
    -- CP-element group 683: successors 
    -- CP-element group 683: marked-successors 
    -- CP-element group 683: 	504 
    -- CP-element group 683: 	516 
    -- CP-element group 683: 	678 
    -- CP-element group 683: 	681 
    -- CP-element group 683:  members (3) 
      -- CP-element group 683: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_sample_completed_
      -- CP-element group 683: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/$exit
      -- CP-element group 683: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/ack
      -- 
    ack_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 683_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1331_inst_ack_0, ack => concat_CP_34_elements(683)); -- 
    -- CP-element group 684:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 684: predecessors 
    -- CP-element group 684: 	682 
    -- CP-element group 684: successors 
    -- CP-element group 684: 	691 
    -- CP-element group 684: marked-successors 
    -- CP-element group 684: 	404 
    -- CP-element group 684: 	682 
    -- CP-element group 684:  members (3) 
      -- CP-element group 684: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_update_completed_
      -- CP-element group 684: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/$exit
      -- CP-element group 684: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/ack
      -- 
    ack_2919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 684_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1331_inst_ack_1, ack => concat_CP_34_elements(684)); -- 
    -- CP-element group 685:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 685: predecessors 
    -- CP-element group 685: 	616 
    -- CP-element group 685: 	624 
    -- CP-element group 685: 	628 
    -- CP-element group 685: 	648 
    -- CP-element group 685: 	652 
    -- CP-element group 685: 	660 
    -- CP-element group 685: marked-predecessors 
    -- CP-element group 685: 	687 
    -- CP-element group 685: successors 
    -- CP-element group 685: 	687 
    -- CP-element group 685:  members (3) 
      -- CP-element group 685: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_sample_start_
      -- CP-element group 685: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/$entry
      -- CP-element group 685: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/rr
      -- 
    rr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(685), ack => type_cast_1346_inst_req_0); -- 
    concat_cp_element_group_685: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_685"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= concat_CP_34_elements(616) & concat_CP_34_elements(624) & concat_CP_34_elements(628) & concat_CP_34_elements(648) & concat_CP_34_elements(652) & concat_CP_34_elements(660) & concat_CP_34_elements(687);
      gj_concat_cp_element_group_685 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(685), clk => clk, reset => reset); --
    end block;
    -- CP-element group 686:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 686: predecessors 
    -- CP-element group 686: marked-predecessors 
    -- CP-element group 686: 	688 
    -- CP-element group 686: successors 
    -- CP-element group 686: 	688 
    -- CP-element group 686:  members (3) 
      -- CP-element group 686: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_update_start_
      -- CP-element group 686: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/$entry
      -- CP-element group 686: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/cr
      -- 
    cr_2932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(686), ack => type_cast_1346_inst_req_1); -- 
    concat_cp_element_group_686: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_686"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(688);
      gj_concat_cp_element_group_686 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(686), clk => clk, reset => reset); --
    end block;
    -- CP-element group 687:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 687: predecessors 
    -- CP-element group 687: 	685 
    -- CP-element group 687: successors 
    -- CP-element group 687: marked-successors 
    -- CP-element group 687: 	614 
    -- CP-element group 687: 	622 
    -- CP-element group 687: 	626 
    -- CP-element group 687: 	646 
    -- CP-element group 687: 	650 
    -- CP-element group 687: 	658 
    -- CP-element group 687: 	685 
    -- CP-element group 687:  members (3) 
      -- CP-element group 687: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_sample_completed_
      -- CP-element group 687: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/$exit
      -- CP-element group 687: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/ra
      -- 
    ra_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 687_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_0, ack => concat_CP_34_elements(687)); -- 
    -- CP-element group 688:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 688: predecessors 
    -- CP-element group 688: 	686 
    -- CP-element group 688: successors 
    -- CP-element group 688: 	317 
    -- CP-element group 688: marked-successors 
    -- CP-element group 688: 	686 
    -- CP-element group 688:  members (3) 
      -- CP-element group 688: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_update_completed_
      -- CP-element group 688: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/$exit
      -- CP-element group 688: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/ca
      -- 
    ca_2933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 688_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_1, ack => concat_CP_34_elements(688)); -- 
    -- CP-element group 689:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 689: predecessors 
    -- CP-element group 689: 	316 
    -- CP-element group 689: successors 
    -- CP-element group 689: 	317 
    -- CP-element group 689:  members (1) 
      -- CP-element group 689: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group concat_CP_34_elements(689) is a control-delay.
    cp_element_689_delay: control_delay_element  generic map(name => " 689_delay", delay_value => 1)  port map(req => concat_CP_34_elements(316), ack => concat_CP_34_elements(689), clk => clk, reset =>reset);
    -- CP-element group 690:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 690: predecessors 
    -- CP-element group 690: 	477 
    -- CP-element group 690: successors 
    -- CP-element group 690: 	585 
    -- CP-element group 690:  members (1) 
      -- CP-element group 690: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_ptr_deref_1113_delay
      -- 
    -- Element group concat_CP_34_elements(690) is a control-delay.
    cp_element_690_delay: control_delay_element  generic map(name => " 690_delay", delay_value => 1)  port map(req => concat_CP_34_elements(477), ack => concat_CP_34_elements(690), clk => clk, reset =>reset);
    -- CP-element group 691:  join  transition  bypass  pipeline-parent 
    -- CP-element group 691: predecessors 
    -- CP-element group 691: 	440 
    -- CP-element group 691: 	463 
    -- CP-element group 691: 	470 
    -- CP-element group 691: 	478 
    -- CP-element group 691: 	486 
    -- CP-element group 691: 	498 
    -- CP-element group 691: 	510 
    -- CP-element group 691: 	530 
    -- CP-element group 691: 	550 
    -- CP-element group 691: 	573 
    -- CP-element group 691: 	580 
    -- CP-element group 691: 	587 
    -- CP-element group 691: 	588 
    -- CP-element group 691: 	620 
    -- CP-element group 691: 	632 
    -- CP-element group 691: 	636 
    -- CP-element group 691: 	644 
    -- CP-element group 691: 	664 
    -- CP-element group 691: 	672 
    -- CP-element group 691: 	676 
    -- CP-element group 691: 	684 
    -- CP-element group 691: successors 
    -- CP-element group 691: 	313 
    -- CP-element group 691:  members (1) 
      -- CP-element group 691: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/$exit
      -- 
    concat_cp_element_group_691: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_691"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= concat_CP_34_elements(440) & concat_CP_34_elements(463) & concat_CP_34_elements(470) & concat_CP_34_elements(478) & concat_CP_34_elements(486) & concat_CP_34_elements(498) & concat_CP_34_elements(510) & concat_CP_34_elements(530) & concat_CP_34_elements(550) & concat_CP_34_elements(573) & concat_CP_34_elements(580) & concat_CP_34_elements(587) & concat_CP_34_elements(588) & concat_CP_34_elements(620) & concat_CP_34_elements(632) & concat_CP_34_elements(636) & concat_CP_34_elements(644) & concat_CP_34_elements(664) & concat_CP_34_elements(672) & concat_CP_34_elements(676) & concat_CP_34_elements(684);
      gj_concat_cp_element_group_691 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(691), clk => clk, reset => reset); --
    end block;
    -- CP-element group 692:  transition  input  bypass  pipeline-parent 
    -- CP-element group 692: predecessors 
    -- CP-element group 692: 	312 
    -- CP-element group 692: successors 
    -- CP-element group 692:  members (2) 
      -- CP-element group 692: 	 branch_block_stmt_23/do_while_stmt_817/loop_exit/$exit
      -- CP-element group 692: 	 branch_block_stmt_23/do_while_stmt_817/loop_exit/ack
      -- 
    ack_2940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 692_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_817_branch_ack_0, ack => concat_CP_34_elements(692)); -- 
    -- CP-element group 693:  transition  input  bypass  pipeline-parent 
    -- CP-element group 693: predecessors 
    -- CP-element group 693: 	312 
    -- CP-element group 693: successors 
    -- CP-element group 693:  members (2) 
      -- CP-element group 693: 	 branch_block_stmt_23/do_while_stmt_817/loop_taken/$exit
      -- CP-element group 693: 	 branch_block_stmt_23/do_while_stmt_817/loop_taken/ack
      -- 
    ack_2944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 693_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_817_branch_ack_1, ack => concat_CP_34_elements(693)); -- 
    -- CP-element group 694:  transition  bypass  pipeline-parent 
    -- CP-element group 694: predecessors 
    -- CP-element group 694: 	310 
    -- CP-element group 694: successors 
    -- CP-element group 694: 	3 
    -- CP-element group 694:  members (1) 
      -- CP-element group 694: 	 branch_block_stmt_23/do_while_stmt_817/$exit
      -- 
    concat_CP_34_elements(694) <= concat_CP_34_elements(310);
    -- CP-element group 695:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 695: predecessors 
    -- CP-element group 695: 	3 
    -- CP-element group 695: successors 
    -- CP-element group 695: 	697 
    -- CP-element group 695: 	698 
    -- CP-element group 695:  members (18) 
      -- CP-element group 695: 	 branch_block_stmt_23/merge_stmt_1363__exit__
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369__entry__
      -- CP-element group 695: 	 branch_block_stmt_23/if_stmt_1359_if_link/$exit
      -- CP-element group 695: 	 branch_block_stmt_23/if_stmt_1359_if_link/if_choice_transition
      -- CP-element group 695: 	 branch_block_stmt_23/ifx_xend297_whilex_xend
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369/$entry
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_sample_start_
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_update_start_
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/$entry
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/rr
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/$entry
      -- CP-element group 695: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/cr
      -- CP-element group 695: 	 branch_block_stmt_23/ifx_xend297_whilex_xend_PhiReq/$entry
      -- CP-element group 695: 	 branch_block_stmt_23/ifx_xend297_whilex_xend_PhiReq/$exit
      -- CP-element group 695: 	 branch_block_stmt_23/merge_stmt_1363_PhiReqMerge
      -- CP-element group 695: 	 branch_block_stmt_23/merge_stmt_1363_PhiAck/$entry
      -- CP-element group 695: 	 branch_block_stmt_23/merge_stmt_1363_PhiAck/$exit
      -- CP-element group 695: 	 branch_block_stmt_23/merge_stmt_1363_PhiAck/dummy
      -- 
    if_choice_transition_2958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 695_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1359_branch_ack_1, ack => concat_CP_34_elements(695)); -- 
    rr_2974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(695), ack => type_cast_1368_inst_req_0); -- 
    cr_2979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(695), ack => type_cast_1368_inst_req_1); -- 
    -- CP-element group 696:  merge  transition  place  input  bypass 
    -- CP-element group 696: predecessors 
    -- CP-element group 696: 	3 
    -- CP-element group 696: successors 
    -- CP-element group 696:  members (5) 
      -- CP-element group 696: 	 branch_block_stmt_23/if_stmt_1359__exit__
      -- CP-element group 696: 	 branch_block_stmt_23/merge_stmt_1363__entry__
      -- CP-element group 696: 	 branch_block_stmt_23/if_stmt_1359_else_link/$exit
      -- CP-element group 696: 	 branch_block_stmt_23/if_stmt_1359_else_link/else_choice_transition
      -- CP-element group 696: 	 branch_block_stmt_23/merge_stmt_1363_dead_link/$entry
      -- 
    else_choice_transition_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 696_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1359_branch_ack_0, ack => concat_CP_34_elements(696)); -- 
    -- CP-element group 697:  transition  input  bypass 
    -- CP-element group 697: predecessors 
    -- CP-element group 697: 	695 
    -- CP-element group 697: successors 
    -- CP-element group 697:  members (3) 
      -- CP-element group 697: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_sample_completed_
      -- CP-element group 697: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/$exit
      -- CP-element group 697: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/ra
      -- 
    ra_2975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 697_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_0, ack => concat_CP_34_elements(697)); -- 
    -- CP-element group 698:  fork  transition  place  input  output  bypass 
    -- CP-element group 698: predecessors 
    -- CP-element group 698: 	695 
    -- CP-element group 698: successors 
    -- CP-element group 698: 	699 
    -- CP-element group 698: 	700 
    -- CP-element group 698: 	702 
    -- CP-element group 698: 	704 
    -- CP-element group 698: 	706 
    -- CP-element group 698: 	708 
    -- CP-element group 698: 	710 
    -- CP-element group 698: 	712 
    -- CP-element group 698: 	714 
    -- CP-element group 698: 	716 
    -- CP-element group 698: 	718 
    -- CP-element group 698:  members (40) 
      -- CP-element group 698: 	 branch_block_stmt_23/assign_stmt_1369__exit__
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480__entry__
      -- CP-element group 698: 	 branch_block_stmt_23/assign_stmt_1369/$exit
      -- CP-element group 698: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_update_completed_
      -- CP-element group 698: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/$exit
      -- CP-element group 698: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/ca
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_sample_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/crr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/ccr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/cr
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_update_start_
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/$entry
      -- CP-element group 698: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/cr
      -- 
    ca_2980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 698_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_1, ack => concat_CP_34_elements(698)); -- 
    crr_2991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => call_stmt_1372_call_req_0); -- 
    ccr_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => call_stmt_1372_call_req_1); -- 
    cr_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1376_inst_req_1); -- 
    cr_3024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1385_inst_req_1); -- 
    cr_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1395_inst_req_1); -- 
    cr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1405_inst_req_1); -- 
    cr_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1415_inst_req_1); -- 
    cr_3080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1425_inst_req_1); -- 
    cr_3094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1435_inst_req_1); -- 
    cr_3108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1445_inst_req_1); -- 
    cr_3122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(698), ack => type_cast_1455_inst_req_1); -- 
    -- CP-element group 699:  transition  input  bypass 
    -- CP-element group 699: predecessors 
    -- CP-element group 699: 	698 
    -- CP-element group 699: successors 
    -- CP-element group 699:  members (3) 
      -- CP-element group 699: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_sample_completed_
      -- CP-element group 699: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/$exit
      -- CP-element group 699: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/cra
      -- 
    cra_2992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 699_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1372_call_ack_0, ack => concat_CP_34_elements(699)); -- 
    -- CP-element group 700:  transition  input  output  bypass 
    -- CP-element group 700: predecessors 
    -- CP-element group 700: 	698 
    -- CP-element group 700: successors 
    -- CP-element group 700: 	701 
    -- CP-element group 700:  members (6) 
      -- CP-element group 700: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_update_completed_
      -- CP-element group 700: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/$exit
      -- CP-element group 700: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/cca
      -- CP-element group 700: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_sample_start_
      -- CP-element group 700: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/$entry
      -- CP-element group 700: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/rr
      -- 
    cca_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 700_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1372_call_ack_1, ack => concat_CP_34_elements(700)); -- 
    rr_3005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(700), ack => type_cast_1376_inst_req_0); -- 
    -- CP-element group 701:  transition  input  bypass 
    -- CP-element group 701: predecessors 
    -- CP-element group 701: 	700 
    -- CP-element group 701: successors 
    -- CP-element group 701:  members (3) 
      -- CP-element group 701: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_sample_completed_
      -- CP-element group 701: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/$exit
      -- CP-element group 701: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/ra
      -- 
    ra_3006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 701_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_0, ack => concat_CP_34_elements(701)); -- 
    -- CP-element group 702:  fork  transition  input  output  bypass 
    -- CP-element group 702: predecessors 
    -- CP-element group 702: 	698 
    -- CP-element group 702: successors 
    -- CP-element group 702: 	703 
    -- CP-element group 702: 	705 
    -- CP-element group 702: 	707 
    -- CP-element group 702: 	709 
    -- CP-element group 702: 	711 
    -- CP-element group 702: 	713 
    -- CP-element group 702: 	715 
    -- CP-element group 702: 	717 
    -- CP-element group 702:  members (27) 
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_update_completed_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/$exit
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/ca
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/rr
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/rr
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/rr
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/rr
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/rr
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/rr
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/rr
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/rr
      -- 
    ca_3011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 702_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_1, ack => concat_CP_34_elements(702)); -- 
    rr_3019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1385_inst_req_0); -- 
    rr_3033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1395_inst_req_0); -- 
    rr_3047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1405_inst_req_0); -- 
    rr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1415_inst_req_0); -- 
    rr_3075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1425_inst_req_0); -- 
    rr_3089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1435_inst_req_0); -- 
    rr_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1445_inst_req_0); -- 
    rr_3117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(702), ack => type_cast_1455_inst_req_0); -- 
    -- CP-element group 703:  transition  input  bypass 
    -- CP-element group 703: predecessors 
    -- CP-element group 703: 	702 
    -- CP-element group 703: successors 
    -- CP-element group 703:  members (3) 
      -- CP-element group 703: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_sample_completed_
      -- CP-element group 703: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/$exit
      -- CP-element group 703: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/ra
      -- 
    ra_3020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 703_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_0, ack => concat_CP_34_elements(703)); -- 
    -- CP-element group 704:  transition  input  bypass 
    -- CP-element group 704: predecessors 
    -- CP-element group 704: 	698 
    -- CP-element group 704: successors 
    -- CP-element group 704: 	739 
    -- CP-element group 704:  members (3) 
      -- CP-element group 704: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_update_completed_
      -- CP-element group 704: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/$exit
      -- CP-element group 704: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/ca
      -- 
    ca_3025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 704_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_1, ack => concat_CP_34_elements(704)); -- 
    -- CP-element group 705:  transition  input  bypass 
    -- CP-element group 705: predecessors 
    -- CP-element group 705: 	702 
    -- CP-element group 705: successors 
    -- CP-element group 705:  members (3) 
      -- CP-element group 705: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_sample_completed_
      -- CP-element group 705: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/$exit
      -- CP-element group 705: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/ra
      -- 
    ra_3034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 705_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_0, ack => concat_CP_34_elements(705)); -- 
    -- CP-element group 706:  transition  input  bypass 
    -- CP-element group 706: predecessors 
    -- CP-element group 706: 	698 
    -- CP-element group 706: successors 
    -- CP-element group 706: 	736 
    -- CP-element group 706:  members (3) 
      -- CP-element group 706: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_update_completed_
      -- CP-element group 706: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/$exit
      -- CP-element group 706: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/ca
      -- 
    ca_3039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 706_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_1, ack => concat_CP_34_elements(706)); -- 
    -- CP-element group 707:  transition  input  bypass 
    -- CP-element group 707: predecessors 
    -- CP-element group 707: 	702 
    -- CP-element group 707: successors 
    -- CP-element group 707:  members (3) 
      -- CP-element group 707: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_sample_completed_
      -- CP-element group 707: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/$exit
      -- CP-element group 707: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/ra
      -- 
    ra_3048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 707_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_0, ack => concat_CP_34_elements(707)); -- 
    -- CP-element group 708:  transition  input  bypass 
    -- CP-element group 708: predecessors 
    -- CP-element group 708: 	698 
    -- CP-element group 708: successors 
    -- CP-element group 708: 	733 
    -- CP-element group 708:  members (3) 
      -- CP-element group 708: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_update_completed_
      -- CP-element group 708: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/$exit
      -- CP-element group 708: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/ca
      -- 
    ca_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 708_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_1, ack => concat_CP_34_elements(708)); -- 
    -- CP-element group 709:  transition  input  bypass 
    -- CP-element group 709: predecessors 
    -- CP-element group 709: 	702 
    -- CP-element group 709: successors 
    -- CP-element group 709:  members (3) 
      -- CP-element group 709: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_sample_completed_
      -- CP-element group 709: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/$exit
      -- CP-element group 709: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/ra
      -- 
    ra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 709_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_0, ack => concat_CP_34_elements(709)); -- 
    -- CP-element group 710:  transition  input  bypass 
    -- CP-element group 710: predecessors 
    -- CP-element group 710: 	698 
    -- CP-element group 710: successors 
    -- CP-element group 710: 	730 
    -- CP-element group 710:  members (3) 
      -- CP-element group 710: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_update_completed_
      -- CP-element group 710: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/$exit
      -- CP-element group 710: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/ca
      -- 
    ca_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 710_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_1, ack => concat_CP_34_elements(710)); -- 
    -- CP-element group 711:  transition  input  bypass 
    -- CP-element group 711: predecessors 
    -- CP-element group 711: 	702 
    -- CP-element group 711: successors 
    -- CP-element group 711:  members (3) 
      -- CP-element group 711: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_sample_completed_
      -- CP-element group 711: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/$exit
      -- CP-element group 711: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/ra
      -- 
    ra_3076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 711_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_0, ack => concat_CP_34_elements(711)); -- 
    -- CP-element group 712:  transition  input  bypass 
    -- CP-element group 712: predecessors 
    -- CP-element group 712: 	698 
    -- CP-element group 712: successors 
    -- CP-element group 712: 	727 
    -- CP-element group 712:  members (3) 
      -- CP-element group 712: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_update_completed_
      -- CP-element group 712: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/$exit
      -- CP-element group 712: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/ca
      -- 
    ca_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 712_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_1, ack => concat_CP_34_elements(712)); -- 
    -- CP-element group 713:  transition  input  bypass 
    -- CP-element group 713: predecessors 
    -- CP-element group 713: 	702 
    -- CP-element group 713: successors 
    -- CP-element group 713:  members (3) 
      -- CP-element group 713: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_sample_completed_
      -- CP-element group 713: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/$exit
      -- CP-element group 713: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/ra
      -- 
    ra_3090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 713_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_0, ack => concat_CP_34_elements(713)); -- 
    -- CP-element group 714:  transition  input  bypass 
    -- CP-element group 714: predecessors 
    -- CP-element group 714: 	698 
    -- CP-element group 714: successors 
    -- CP-element group 714: 	724 
    -- CP-element group 714:  members (3) 
      -- CP-element group 714: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_update_completed_
      -- CP-element group 714: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/$exit
      -- CP-element group 714: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/ca
      -- 
    ca_3095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 714_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_1, ack => concat_CP_34_elements(714)); -- 
    -- CP-element group 715:  transition  input  bypass 
    -- CP-element group 715: predecessors 
    -- CP-element group 715: 	702 
    -- CP-element group 715: successors 
    -- CP-element group 715:  members (3) 
      -- CP-element group 715: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_sample_completed_
      -- CP-element group 715: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/$exit
      -- CP-element group 715: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/ra
      -- 
    ra_3104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 715_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_0, ack => concat_CP_34_elements(715)); -- 
    -- CP-element group 716:  transition  input  bypass 
    -- CP-element group 716: predecessors 
    -- CP-element group 716: 	698 
    -- CP-element group 716: successors 
    -- CP-element group 716: 	721 
    -- CP-element group 716:  members (3) 
      -- CP-element group 716: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_update_completed_
      -- CP-element group 716: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/$exit
      -- CP-element group 716: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/ca
      -- 
    ca_3109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 716_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_1, ack => concat_CP_34_elements(716)); -- 
    -- CP-element group 717:  transition  input  bypass 
    -- CP-element group 717: predecessors 
    -- CP-element group 717: 	702 
    -- CP-element group 717: successors 
    -- CP-element group 717:  members (3) 
      -- CP-element group 717: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_sample_completed_
      -- CP-element group 717: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/$exit
      -- CP-element group 717: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/ra
      -- 
    ra_3118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 717_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_0, ack => concat_CP_34_elements(717)); -- 
    -- CP-element group 718:  transition  input  output  bypass 
    -- CP-element group 718: predecessors 
    -- CP-element group 718: 	698 
    -- CP-element group 718: successors 
    -- CP-element group 718: 	719 
    -- CP-element group 718:  members (6) 
      -- CP-element group 718: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_update_completed_
      -- CP-element group 718: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/$exit
      -- CP-element group 718: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/ca
      -- CP-element group 718: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_sample_start_
      -- CP-element group 718: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/$entry
      -- CP-element group 718: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/req
      -- 
    ca_3123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 718_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_1, ack => concat_CP_34_elements(718)); -- 
    req_3131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(718), ack => WPIPE_Concat_output_pipe_1457_inst_req_0); -- 
    -- CP-element group 719:  transition  input  output  bypass 
    -- CP-element group 719: predecessors 
    -- CP-element group 719: 	718 
    -- CP-element group 719: successors 
    -- CP-element group 719: 	720 
    -- CP-element group 719:  members (6) 
      -- CP-element group 719: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/req
      -- CP-element group 719: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/$entry
      -- CP-element group 719: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_sample_completed_
      -- CP-element group 719: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_update_start_
      -- CP-element group 719: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/$exit
      -- CP-element group 719: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/ack
      -- 
    ack_3132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 719_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1457_inst_ack_0, ack => concat_CP_34_elements(719)); -- 
    req_3136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(719), ack => WPIPE_Concat_output_pipe_1457_inst_req_1); -- 
    -- CP-element group 720:  transition  input  bypass 
    -- CP-element group 720: predecessors 
    -- CP-element group 720: 	719 
    -- CP-element group 720: successors 
    -- CP-element group 720: 	721 
    -- CP-element group 720:  members (3) 
      -- CP-element group 720: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/ack
      -- CP-element group 720: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/$exit
      -- CP-element group 720: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_update_completed_
      -- 
    ack_3137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 720_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1457_inst_ack_1, ack => concat_CP_34_elements(720)); -- 
    -- CP-element group 721:  join  transition  output  bypass 
    -- CP-element group 721: predecessors 
    -- CP-element group 721: 	716 
    -- CP-element group 721: 	720 
    -- CP-element group 721: successors 
    -- CP-element group 721: 	722 
    -- CP-element group 721:  members (3) 
      -- CP-element group 721: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/req
      -- CP-element group 721: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/$entry
      -- CP-element group 721: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_sample_start_
      -- 
    req_3145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(721), ack => WPIPE_Concat_output_pipe_1460_inst_req_0); -- 
    concat_cp_element_group_721: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_721"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(716) & concat_CP_34_elements(720);
      gj_concat_cp_element_group_721 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(721), clk => clk, reset => reset); --
    end block;
    -- CP-element group 722:  transition  input  output  bypass 
    -- CP-element group 722: predecessors 
    -- CP-element group 722: 	721 
    -- CP-element group 722: successors 
    -- CP-element group 722: 	723 
    -- CP-element group 722:  members (6) 
      -- CP-element group 722: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/req
      -- CP-element group 722: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/ack
      -- CP-element group 722: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/$exit
      -- CP-element group 722: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_update_start_
      -- CP-element group 722: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_sample_completed_
      -- 
    ack_3146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 722_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1460_inst_ack_0, ack => concat_CP_34_elements(722)); -- 
    req_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(722), ack => WPIPE_Concat_output_pipe_1460_inst_req_1); -- 
    -- CP-element group 723:  transition  input  bypass 
    -- CP-element group 723: predecessors 
    -- CP-element group 723: 	722 
    -- CP-element group 723: successors 
    -- CP-element group 723: 	724 
    -- CP-element group 723:  members (3) 
      -- CP-element group 723: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/$exit
      -- CP-element group 723: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/ack
      -- CP-element group 723: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_update_completed_
      -- 
    ack_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 723_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1460_inst_ack_1, ack => concat_CP_34_elements(723)); -- 
    -- CP-element group 724:  join  transition  output  bypass 
    -- CP-element group 724: predecessors 
    -- CP-element group 724: 	714 
    -- CP-element group 724: 	723 
    -- CP-element group 724: successors 
    -- CP-element group 724: 	725 
    -- CP-element group 724:  members (3) 
      -- CP-element group 724: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_sample_start_
      -- CP-element group 724: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/$entry
      -- CP-element group 724: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/req
      -- 
    req_3159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(724), ack => WPIPE_Concat_output_pipe_1463_inst_req_0); -- 
    concat_cp_element_group_724: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_724"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(714) & concat_CP_34_elements(723);
      gj_concat_cp_element_group_724 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(724), clk => clk, reset => reset); --
    end block;
    -- CP-element group 725:  transition  input  output  bypass 
    -- CP-element group 725: predecessors 
    -- CP-element group 725: 	724 
    -- CP-element group 725: successors 
    -- CP-element group 725: 	726 
    -- CP-element group 725:  members (6) 
      -- CP-element group 725: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_sample_completed_
      -- CP-element group 725: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_update_start_
      -- CP-element group 725: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/$exit
      -- CP-element group 725: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/ack
      -- CP-element group 725: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/$entry
      -- CP-element group 725: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/req
      -- 
    ack_3160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 725_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1463_inst_ack_0, ack => concat_CP_34_elements(725)); -- 
    req_3164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(725), ack => WPIPE_Concat_output_pipe_1463_inst_req_1); -- 
    -- CP-element group 726:  transition  input  bypass 
    -- CP-element group 726: predecessors 
    -- CP-element group 726: 	725 
    -- CP-element group 726: successors 
    -- CP-element group 726: 	727 
    -- CP-element group 726:  members (3) 
      -- CP-element group 726: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_update_completed_
      -- CP-element group 726: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/$exit
      -- CP-element group 726: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/ack
      -- 
    ack_3165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 726_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1463_inst_ack_1, ack => concat_CP_34_elements(726)); -- 
    -- CP-element group 727:  join  transition  output  bypass 
    -- CP-element group 727: predecessors 
    -- CP-element group 727: 	712 
    -- CP-element group 727: 	726 
    -- CP-element group 727: successors 
    -- CP-element group 727: 	728 
    -- CP-element group 727:  members (3) 
      -- CP-element group 727: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_sample_start_
      -- CP-element group 727: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/$entry
      -- CP-element group 727: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/req
      -- 
    req_3173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(727), ack => WPIPE_Concat_output_pipe_1466_inst_req_0); -- 
    concat_cp_element_group_727: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_727"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(712) & concat_CP_34_elements(726);
      gj_concat_cp_element_group_727 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(727), clk => clk, reset => reset); --
    end block;
    -- CP-element group 728:  transition  input  output  bypass 
    -- CP-element group 728: predecessors 
    -- CP-element group 728: 	727 
    -- CP-element group 728: successors 
    -- CP-element group 728: 	729 
    -- CP-element group 728:  members (6) 
      -- CP-element group 728: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_sample_completed_
      -- CP-element group 728: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_update_start_
      -- CP-element group 728: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/$exit
      -- CP-element group 728: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/ack
      -- CP-element group 728: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/$entry
      -- CP-element group 728: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/req
      -- 
    ack_3174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 728_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1466_inst_ack_0, ack => concat_CP_34_elements(728)); -- 
    req_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(728), ack => WPIPE_Concat_output_pipe_1466_inst_req_1); -- 
    -- CP-element group 729:  transition  input  bypass 
    -- CP-element group 729: predecessors 
    -- CP-element group 729: 	728 
    -- CP-element group 729: successors 
    -- CP-element group 729: 	730 
    -- CP-element group 729:  members (3) 
      -- CP-element group 729: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_update_completed_
      -- CP-element group 729: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/$exit
      -- CP-element group 729: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/ack
      -- 
    ack_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 729_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1466_inst_ack_1, ack => concat_CP_34_elements(729)); -- 
    -- CP-element group 730:  join  transition  output  bypass 
    -- CP-element group 730: predecessors 
    -- CP-element group 730: 	710 
    -- CP-element group 730: 	729 
    -- CP-element group 730: successors 
    -- CP-element group 730: 	731 
    -- CP-element group 730:  members (3) 
      -- CP-element group 730: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/$entry
      -- CP-element group 730: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/req
      -- CP-element group 730: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_sample_start_
      -- 
    req_3187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(730), ack => WPIPE_Concat_output_pipe_1469_inst_req_0); -- 
    concat_cp_element_group_730: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_730"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(710) & concat_CP_34_elements(729);
      gj_concat_cp_element_group_730 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(730), clk => clk, reset => reset); --
    end block;
    -- CP-element group 731:  transition  input  output  bypass 
    -- CP-element group 731: predecessors 
    -- CP-element group 731: 	730 
    -- CP-element group 731: successors 
    -- CP-element group 731: 	732 
    -- CP-element group 731:  members (6) 
      -- CP-element group 731: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_sample_completed_
      -- CP-element group 731: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_update_start_
      -- CP-element group 731: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/$exit
      -- CP-element group 731: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/ack
      -- CP-element group 731: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/$entry
      -- CP-element group 731: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/req
      -- 
    ack_3188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 731_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1469_inst_ack_0, ack => concat_CP_34_elements(731)); -- 
    req_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(731), ack => WPIPE_Concat_output_pipe_1469_inst_req_1); -- 
    -- CP-element group 732:  transition  input  bypass 
    -- CP-element group 732: predecessors 
    -- CP-element group 732: 	731 
    -- CP-element group 732: successors 
    -- CP-element group 732: 	733 
    -- CP-element group 732:  members (3) 
      -- CP-element group 732: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_update_completed_
      -- CP-element group 732: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/ack
      -- CP-element group 732: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/$exit
      -- 
    ack_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 732_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1469_inst_ack_1, ack => concat_CP_34_elements(732)); -- 
    -- CP-element group 733:  join  transition  output  bypass 
    -- CP-element group 733: predecessors 
    -- CP-element group 733: 	708 
    -- CP-element group 733: 	732 
    -- CP-element group 733: successors 
    -- CP-element group 733: 	734 
    -- CP-element group 733:  members (3) 
      -- CP-element group 733: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/$entry
      -- CP-element group 733: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/req
      -- CP-element group 733: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_sample_start_
      -- 
    req_3201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(733), ack => WPIPE_Concat_output_pipe_1472_inst_req_0); -- 
    concat_cp_element_group_733: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_733"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(708) & concat_CP_34_elements(732);
      gj_concat_cp_element_group_733 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(733), clk => clk, reset => reset); --
    end block;
    -- CP-element group 734:  transition  input  output  bypass 
    -- CP-element group 734: predecessors 
    -- CP-element group 734: 	733 
    -- CP-element group 734: successors 
    -- CP-element group 734: 	735 
    -- CP-element group 734:  members (6) 
      -- CP-element group 734: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/$exit
      -- CP-element group 734: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/ack
      -- CP-element group 734: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/$entry
      -- CP-element group 734: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/req
      -- CP-element group 734: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_update_start_
      -- CP-element group 734: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_sample_completed_
      -- 
    ack_3202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 734_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1472_inst_ack_0, ack => concat_CP_34_elements(734)); -- 
    req_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(734), ack => WPIPE_Concat_output_pipe_1472_inst_req_1); -- 
    -- CP-element group 735:  transition  input  bypass 
    -- CP-element group 735: predecessors 
    -- CP-element group 735: 	734 
    -- CP-element group 735: successors 
    -- CP-element group 735: 	736 
    -- CP-element group 735:  members (3) 
      -- CP-element group 735: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/$exit
      -- CP-element group 735: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/ack
      -- CP-element group 735: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_update_completed_
      -- 
    ack_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 735_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1472_inst_ack_1, ack => concat_CP_34_elements(735)); -- 
    -- CP-element group 736:  join  transition  output  bypass 
    -- CP-element group 736: predecessors 
    -- CP-element group 736: 	706 
    -- CP-element group 736: 	735 
    -- CP-element group 736: successors 
    -- CP-element group 736: 	737 
    -- CP-element group 736:  members (3) 
      -- CP-element group 736: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_sample_start_
      -- CP-element group 736: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/$entry
      -- CP-element group 736: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/req
      -- 
    req_3215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(736), ack => WPIPE_Concat_output_pipe_1475_inst_req_0); -- 
    concat_cp_element_group_736: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_736"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(706) & concat_CP_34_elements(735);
      gj_concat_cp_element_group_736 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(736), clk => clk, reset => reset); --
    end block;
    -- CP-element group 737:  transition  input  output  bypass 
    -- CP-element group 737: predecessors 
    -- CP-element group 737: 	736 
    -- CP-element group 737: successors 
    -- CP-element group 737: 	738 
    -- CP-element group 737:  members (6) 
      -- CP-element group 737: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_sample_completed_
      -- CP-element group 737: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_update_start_
      -- CP-element group 737: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/$exit
      -- CP-element group 737: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/ack
      -- CP-element group 737: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/req
      -- 
    ack_3216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 737_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1475_inst_ack_0, ack => concat_CP_34_elements(737)); -- 
    req_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(737), ack => WPIPE_Concat_output_pipe_1475_inst_req_1); -- 
    -- CP-element group 738:  transition  input  bypass 
    -- CP-element group 738: predecessors 
    -- CP-element group 738: 	737 
    -- CP-element group 738: successors 
    -- CP-element group 738: 	739 
    -- CP-element group 738:  members (3) 
      -- CP-element group 738: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_update_completed_
      -- CP-element group 738: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/$exit
      -- CP-element group 738: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/ack
      -- 
    ack_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 738_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1475_inst_ack_1, ack => concat_CP_34_elements(738)); -- 
    -- CP-element group 739:  join  transition  output  bypass 
    -- CP-element group 739: predecessors 
    -- CP-element group 739: 	704 
    -- CP-element group 739: 	738 
    -- CP-element group 739: successors 
    -- CP-element group 739: 	740 
    -- CP-element group 739:  members (3) 
      -- CP-element group 739: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/req
      -- CP-element group 739: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_sample_start_
      -- CP-element group 739: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/$entry
      -- 
    req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(739), ack => WPIPE_Concat_output_pipe_1478_inst_req_0); -- 
    concat_cp_element_group_739: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_739"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(704) & concat_CP_34_elements(738);
      gj_concat_cp_element_group_739 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(739), clk => clk, reset => reset); --
    end block;
    -- CP-element group 740:  transition  input  output  bypass 
    -- CP-element group 740: predecessors 
    -- CP-element group 740: 	739 
    -- CP-element group 740: successors 
    -- CP-element group 740: 	741 
    -- CP-element group 740:  members (6) 
      -- CP-element group 740: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/ack
      -- CP-element group 740: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/$entry
      -- CP-element group 740: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/req
      -- CP-element group 740: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_sample_completed_
      -- CP-element group 740: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_update_start_
      -- CP-element group 740: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/$exit
      -- 
    ack_3230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 740_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1478_inst_ack_0, ack => concat_CP_34_elements(740)); -- 
    req_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(740), ack => WPIPE_Concat_output_pipe_1478_inst_req_1); -- 
    -- CP-element group 741:  branch  transition  place  input  output  bypass 
    -- CP-element group 741: predecessors 
    -- CP-element group 741: 	740 
    -- CP-element group 741: successors 
    -- CP-element group 741: 	742 
    -- CP-element group 741: 	743 
    -- CP-element group 741:  members (17) 
      -- CP-element group 741: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480__exit__
      -- CP-element group 741: 	 branch_block_stmt_23/assign_stmt_1487__entry__
      -- CP-element group 741: 	 branch_block_stmt_23/assign_stmt_1487__exit__
      -- CP-element group 741: 	 branch_block_stmt_23/if_stmt_1488__entry__
      -- CP-element group 741: 	 branch_block_stmt_23/R_cmp378460_1489_place
      -- CP-element group 741: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/$exit
      -- CP-element group 741: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/ack
      -- CP-element group 741: 	 branch_block_stmt_23/assign_stmt_1487/$entry
      -- CP-element group 741: 	 branch_block_stmt_23/assign_stmt_1487/$exit
      -- CP-element group 741: 	 branch_block_stmt_23/if_stmt_1488_dead_link/$entry
      -- CP-element group 741: 	 branch_block_stmt_23/if_stmt_1488_eval_test/$entry
      -- CP-element group 741: 	 branch_block_stmt_23/if_stmt_1488_eval_test/$exit
      -- CP-element group 741: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_update_completed_
      -- CP-element group 741: 	 branch_block_stmt_23/if_stmt_1488_else_link/$entry
      -- CP-element group 741: 	 branch_block_stmt_23/if_stmt_1488_if_link/$entry
      -- CP-element group 741: 	 branch_block_stmt_23/if_stmt_1488_eval_test/branch_req
      -- CP-element group 741: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/$exit
      -- 
    ack_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 741_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1478_inst_ack_1, ack => concat_CP_34_elements(741)); -- 
    branch_req_3246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(741), ack => if_stmt_1488_branch_req_0); -- 
    -- CP-element group 742:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 742: predecessors 
    -- CP-element group 742: 	741 
    -- CP-element group 742: successors 
    -- CP-element group 742: 	744 
    -- CP-element group 742: 	745 
    -- CP-element group 742:  members (18) 
      -- CP-element group 742: 	 branch_block_stmt_23/merge_stmt_1494__exit__
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523__entry__
      -- CP-element group 742: 	 branch_block_stmt_23/whilex_xend_bbx_xnph
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_update_start_
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/$entry
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/rr
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_sample_start_
      -- CP-element group 742: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/$entry
      -- CP-element group 742: 	 branch_block_stmt_23/if_stmt_1488_if_link/if_choice_transition
      -- CP-element group 742: 	 branch_block_stmt_23/if_stmt_1488_if_link/$exit
      -- CP-element group 742: 	 branch_block_stmt_23/whilex_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 742: 	 branch_block_stmt_23/whilex_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 742: 	 branch_block_stmt_23/merge_stmt_1494_PhiReqMerge
      -- CP-element group 742: 	 branch_block_stmt_23/merge_stmt_1494_PhiAck/$entry
      -- CP-element group 742: 	 branch_block_stmt_23/merge_stmt_1494_PhiAck/$exit
      -- CP-element group 742: 	 branch_block_stmt_23/merge_stmt_1494_PhiAck/dummy
      -- 
    if_choice_transition_3251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 742_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_1, ack => concat_CP_34_elements(742)); -- 
    rr_3268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(742), ack => type_cast_1509_inst_req_0); -- 
    cr_3273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(742), ack => type_cast_1509_inst_req_1); -- 
    -- CP-element group 743:  transition  place  input  bypass 
    -- CP-element group 743: predecessors 
    -- CP-element group 743: 	741 
    -- CP-element group 743: successors 
    -- CP-element group 743: 	802 
    -- CP-element group 743:  members (5) 
      -- CP-element group 743: 	 branch_block_stmt_23/whilex_xend_forx_xend453
      -- CP-element group 743: 	 branch_block_stmt_23/if_stmt_1488_else_link/else_choice_transition
      -- CP-element group 743: 	 branch_block_stmt_23/if_stmt_1488_else_link/$exit
      -- CP-element group 743: 	 branch_block_stmt_23/whilex_xend_forx_xend453_PhiReq/$entry
      -- CP-element group 743: 	 branch_block_stmt_23/whilex_xend_forx_xend453_PhiReq/$exit
      -- 
    else_choice_transition_3255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 743_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_0, ack => concat_CP_34_elements(743)); -- 
    -- CP-element group 744:  transition  input  bypass 
    -- CP-element group 744: predecessors 
    -- CP-element group 744: 	742 
    -- CP-element group 744: successors 
    -- CP-element group 744:  members (3) 
      -- CP-element group 744: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/$exit
      -- CP-element group 744: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/ra
      -- CP-element group 744: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_sample_completed_
      -- 
    ra_3269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 744_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_0, ack => concat_CP_34_elements(744)); -- 
    -- CP-element group 745:  transition  place  input  bypass 
    -- CP-element group 745: predecessors 
    -- CP-element group 745: 	742 
    -- CP-element group 745: successors 
    -- CP-element group 745: 	796 
    -- CP-element group 745:  members (9) 
      -- CP-element group 745: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_update_completed_
      -- CP-element group 745: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523__exit__
      -- CP-element group 745: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380
      -- CP-element group 745: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/$exit
      -- CP-element group 745: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/ca
      -- CP-element group 745: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/$exit
      -- CP-element group 745: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/$entry
      -- CP-element group 745: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/phi_stmt_1526/$entry
      -- CP-element group 745: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$entry
      -- 
    ca_3274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 745_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_1, ack => concat_CP_34_elements(745)); -- 
    -- CP-element group 746:  transition  input  bypass 
    -- CP-element group 746: predecessors 
    -- CP-element group 746: 	801 
    -- CP-element group 746: successors 
    -- CP-element group 746: 	791 
    -- CP-element group 746:  members (3) 
      -- CP-element group 746: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/ack
      -- CP-element group 746: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_sample_complete
      -- CP-element group 746: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/$exit
      -- 
    ack_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 746_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1538_index_offset_ack_0, ack => concat_CP_34_elements(746)); -- 
    -- CP-element group 747:  transition  input  output  bypass 
    -- CP-element group 747: predecessors 
    -- CP-element group 747: 	801 
    -- CP-element group 747: successors 
    -- CP-element group 747: 	748 
    -- CP-element group 747:  members (11) 
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/$exit
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_sample_start_
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/ack
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_root_address_calculated
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/$entry
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_offset_calculated
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/$exit
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/sum_rename_req
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/sum_rename_ack
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/$entry
      -- CP-element group 747: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/req
      -- 
    ack_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 747_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1538_index_offset_ack_1, ack => concat_CP_34_elements(747)); -- 
    req_3317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(747), ack => addr_of_1539_final_reg_req_0); -- 
    -- CP-element group 748:  transition  input  bypass 
    -- CP-element group 748: predecessors 
    -- CP-element group 748: 	747 
    -- CP-element group 748: successors 
    -- CP-element group 748:  members (3) 
      -- CP-element group 748: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_sample_completed_
      -- CP-element group 748: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/$exit
      -- CP-element group 748: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/ack
      -- 
    ack_3318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 748_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1539_final_reg_ack_0, ack => concat_CP_34_elements(748)); -- 
    -- CP-element group 749:  join  fork  transition  input  output  bypass 
    -- CP-element group 749: predecessors 
    -- CP-element group 749: 	801 
    -- CP-element group 749: successors 
    -- CP-element group 749: 	750 
    -- CP-element group 749:  members (24) 
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_address_calculated
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_address_calculated
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_root_address_calculated
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_address_resized
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/$entry
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/$exit
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/base_resize_req
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/base_resize_ack
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/$entry
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_update_completed_
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/$exit
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/sum_rename_req
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/sum_rename_ack
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/$entry
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/$exit
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/root_register_req
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/root_register_ack
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/$entry
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/$entry
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/$entry
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/rr
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_sample_start_
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/ack
      -- CP-element group 749: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/$exit
      -- 
    ack_3323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 749_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1539_final_reg_ack_1, ack => concat_CP_34_elements(749)); -- 
    rr_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(749), ack => ptr_deref_1543_load_0_req_0); -- 
    -- CP-element group 750:  transition  input  bypass 
    -- CP-element group 750: predecessors 
    -- CP-element group 750: 	749 
    -- CP-element group 750: successors 
    -- CP-element group 750:  members (5) 
      -- CP-element group 750: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/$exit
      -- CP-element group 750: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/$exit
      -- CP-element group 750: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/$exit
      -- CP-element group 750: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/ra
      -- CP-element group 750: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_sample_completed_
      -- 
    ra_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 750_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_load_0_ack_0, ack => concat_CP_34_elements(750)); -- 
    -- CP-element group 751:  fork  transition  input  output  bypass 
    -- CP-element group 751: predecessors 
    -- CP-element group 751: 	801 
    -- CP-element group 751: successors 
    -- CP-element group 751: 	752 
    -- CP-element group 751: 	754 
    -- CP-element group 751: 	756 
    -- CP-element group 751: 	758 
    -- CP-element group 751: 	760 
    -- CP-element group 751: 	762 
    -- CP-element group 751: 	764 
    -- CP-element group 751: 	766 
    -- CP-element group 751:  members (33) 
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/ca
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_update_completed_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/$exit
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/merge_req
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/merge_ack
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/rr
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/rr
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/rr
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/rr
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/rr
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/rr
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/$exit
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/$exit
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/$exit
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/rr
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_sample_start_
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/$entry
      -- CP-element group 751: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/rr
      -- 
    ca_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 751_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_load_0_ack_1, ack => concat_CP_34_elements(751)); -- 
    rr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1547_inst_req_0); -- 
    rr_3395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1557_inst_req_0); -- 
    rr_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1567_inst_req_0); -- 
    rr_3423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1577_inst_req_0); -- 
    rr_3437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1587_inst_req_0); -- 
    rr_3451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1597_inst_req_0); -- 
    rr_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1607_inst_req_0); -- 
    rr_3479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(751), ack => type_cast_1617_inst_req_0); -- 
    -- CP-element group 752:  transition  input  bypass 
    -- CP-element group 752: predecessors 
    -- CP-element group 752: 	751 
    -- CP-element group 752: successors 
    -- CP-element group 752:  members (3) 
      -- CP-element group 752: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_sample_completed_
      -- CP-element group 752: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/$exit
      -- CP-element group 752: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/ra
      -- 
    ra_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 752_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1547_inst_ack_0, ack => concat_CP_34_elements(752)); -- 
    -- CP-element group 753:  transition  input  bypass 
    -- CP-element group 753: predecessors 
    -- CP-element group 753: 	801 
    -- CP-element group 753: successors 
    -- CP-element group 753: 	788 
    -- CP-element group 753:  members (3) 
      -- CP-element group 753: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_update_completed_
      -- CP-element group 753: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/$exit
      -- CP-element group 753: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/ca
      -- 
    ca_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 753_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1547_inst_ack_1, ack => concat_CP_34_elements(753)); -- 
    -- CP-element group 754:  transition  input  bypass 
    -- CP-element group 754: predecessors 
    -- CP-element group 754: 	751 
    -- CP-element group 754: successors 
    -- CP-element group 754:  members (3) 
      -- CP-element group 754: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/$exit
      -- CP-element group 754: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_sample_completed_
      -- CP-element group 754: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/ra
      -- 
    ra_3396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 754_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_0, ack => concat_CP_34_elements(754)); -- 
    -- CP-element group 755:  transition  input  bypass 
    -- CP-element group 755: predecessors 
    -- CP-element group 755: 	801 
    -- CP-element group 755: successors 
    -- CP-element group 755: 	785 
    -- CP-element group 755:  members (3) 
      -- CP-element group 755: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_update_completed_
      -- CP-element group 755: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/ca
      -- CP-element group 755: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/$exit
      -- 
    ca_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 755_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_1, ack => concat_CP_34_elements(755)); -- 
    -- CP-element group 756:  transition  input  bypass 
    -- CP-element group 756: predecessors 
    -- CP-element group 756: 	751 
    -- CP-element group 756: successors 
    -- CP-element group 756:  members (3) 
      -- CP-element group 756: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/$exit
      -- CP-element group 756: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/ra
      -- CP-element group 756: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_sample_completed_
      -- 
    ra_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 756_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_0, ack => concat_CP_34_elements(756)); -- 
    -- CP-element group 757:  transition  input  bypass 
    -- CP-element group 757: predecessors 
    -- CP-element group 757: 	801 
    -- CP-element group 757: successors 
    -- CP-element group 757: 	782 
    -- CP-element group 757:  members (3) 
      -- CP-element group 757: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_update_completed_
      -- CP-element group 757: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/$exit
      -- CP-element group 757: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/ca
      -- 
    ca_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 757_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_1, ack => concat_CP_34_elements(757)); -- 
    -- CP-element group 758:  transition  input  bypass 
    -- CP-element group 758: predecessors 
    -- CP-element group 758: 	751 
    -- CP-element group 758: successors 
    -- CP-element group 758:  members (3) 
      -- CP-element group 758: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_sample_completed_
      -- CP-element group 758: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/$exit
      -- CP-element group 758: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/ra
      -- 
    ra_3424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 758_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_0, ack => concat_CP_34_elements(758)); -- 
    -- CP-element group 759:  transition  input  bypass 
    -- CP-element group 759: predecessors 
    -- CP-element group 759: 	801 
    -- CP-element group 759: successors 
    -- CP-element group 759: 	779 
    -- CP-element group 759:  members (3) 
      -- CP-element group 759: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_update_completed_
      -- CP-element group 759: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/ca
      -- CP-element group 759: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/$exit
      -- 
    ca_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 759_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_1, ack => concat_CP_34_elements(759)); -- 
    -- CP-element group 760:  transition  input  bypass 
    -- CP-element group 760: predecessors 
    -- CP-element group 760: 	751 
    -- CP-element group 760: successors 
    -- CP-element group 760:  members (3) 
      -- CP-element group 760: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/$exit
      -- CP-element group 760: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/ra
      -- CP-element group 760: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_sample_completed_
      -- 
    ra_3438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 760_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_0, ack => concat_CP_34_elements(760)); -- 
    -- CP-element group 761:  transition  input  bypass 
    -- CP-element group 761: predecessors 
    -- CP-element group 761: 	801 
    -- CP-element group 761: successors 
    -- CP-element group 761: 	776 
    -- CP-element group 761:  members (3) 
      -- CP-element group 761: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_update_completed_
      -- CP-element group 761: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/$exit
      -- CP-element group 761: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/ca
      -- 
    ca_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 761_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_1, ack => concat_CP_34_elements(761)); -- 
    -- CP-element group 762:  transition  input  bypass 
    -- CP-element group 762: predecessors 
    -- CP-element group 762: 	751 
    -- CP-element group 762: successors 
    -- CP-element group 762:  members (3) 
      -- CP-element group 762: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_sample_completed_
      -- CP-element group 762: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/$exit
      -- CP-element group 762: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/ra
      -- 
    ra_3452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 762_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_0, ack => concat_CP_34_elements(762)); -- 
    -- CP-element group 763:  transition  input  bypass 
    -- CP-element group 763: predecessors 
    -- CP-element group 763: 	801 
    -- CP-element group 763: successors 
    -- CP-element group 763: 	773 
    -- CP-element group 763:  members (3) 
      -- CP-element group 763: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/ca
      -- CP-element group 763: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_update_completed_
      -- CP-element group 763: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/$exit
      -- 
    ca_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 763_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_1, ack => concat_CP_34_elements(763)); -- 
    -- CP-element group 764:  transition  input  bypass 
    -- CP-element group 764: predecessors 
    -- CP-element group 764: 	751 
    -- CP-element group 764: successors 
    -- CP-element group 764:  members (3) 
      -- CP-element group 764: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_sample_completed_
      -- CP-element group 764: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/$exit
      -- CP-element group 764: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/ra
      -- 
    ra_3466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 764_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_0, ack => concat_CP_34_elements(764)); -- 
    -- CP-element group 765:  transition  input  bypass 
    -- CP-element group 765: predecessors 
    -- CP-element group 765: 	801 
    -- CP-element group 765: successors 
    -- CP-element group 765: 	770 
    -- CP-element group 765:  members (3) 
      -- CP-element group 765: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_update_completed_
      -- CP-element group 765: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/$exit
      -- CP-element group 765: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/ca
      -- 
    ca_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 765_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_1, ack => concat_CP_34_elements(765)); -- 
    -- CP-element group 766:  transition  input  bypass 
    -- CP-element group 766: predecessors 
    -- CP-element group 766: 	751 
    -- CP-element group 766: successors 
    -- CP-element group 766:  members (3) 
      -- CP-element group 766: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_sample_completed_
      -- CP-element group 766: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/$exit
      -- CP-element group 766: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/ra
      -- 
    ra_3480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 766_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_0, ack => concat_CP_34_elements(766)); -- 
    -- CP-element group 767:  transition  input  output  bypass 
    -- CP-element group 767: predecessors 
    -- CP-element group 767: 	801 
    -- CP-element group 767: successors 
    -- CP-element group 767: 	768 
    -- CP-element group 767:  members (6) 
      -- CP-element group 767: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_update_completed_
      -- CP-element group 767: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/$exit
      -- CP-element group 767: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/ca
      -- CP-element group 767: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_sample_start_
      -- CP-element group 767: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/$entry
      -- CP-element group 767: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/req
      -- 
    ca_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 767_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_1, ack => concat_CP_34_elements(767)); -- 
    req_3493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(767), ack => WPIPE_Concat_output_pipe_1619_inst_req_0); -- 
    -- CP-element group 768:  transition  input  output  bypass 
    -- CP-element group 768: predecessors 
    -- CP-element group 768: 	767 
    -- CP-element group 768: successors 
    -- CP-element group 768: 	769 
    -- CP-element group 768:  members (6) 
      -- CP-element group 768: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_sample_completed_
      -- CP-element group 768: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_update_start_
      -- CP-element group 768: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/$exit
      -- CP-element group 768: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/ack
      -- CP-element group 768: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/$entry
      -- CP-element group 768: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/req
      -- 
    ack_3494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 768_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1619_inst_ack_0, ack => concat_CP_34_elements(768)); -- 
    req_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(768), ack => WPIPE_Concat_output_pipe_1619_inst_req_1); -- 
    -- CP-element group 769:  transition  input  bypass 
    -- CP-element group 769: predecessors 
    -- CP-element group 769: 	768 
    -- CP-element group 769: successors 
    -- CP-element group 769: 	770 
    -- CP-element group 769:  members (3) 
      -- CP-element group 769: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_update_completed_
      -- CP-element group 769: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/$exit
      -- CP-element group 769: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/ack
      -- 
    ack_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 769_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1619_inst_ack_1, ack => concat_CP_34_elements(769)); -- 
    -- CP-element group 770:  join  transition  output  bypass 
    -- CP-element group 770: predecessors 
    -- CP-element group 770: 	765 
    -- CP-element group 770: 	769 
    -- CP-element group 770: successors 
    -- CP-element group 770: 	771 
    -- CP-element group 770:  members (3) 
      -- CP-element group 770: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_sample_start_
      -- CP-element group 770: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/$entry
      -- CP-element group 770: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/req
      -- 
    req_3507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(770), ack => WPIPE_Concat_output_pipe_1622_inst_req_0); -- 
    concat_cp_element_group_770: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_770"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(765) & concat_CP_34_elements(769);
      gj_concat_cp_element_group_770 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(770), clk => clk, reset => reset); --
    end block;
    -- CP-element group 771:  transition  input  output  bypass 
    -- CP-element group 771: predecessors 
    -- CP-element group 771: 	770 
    -- CP-element group 771: successors 
    -- CP-element group 771: 	772 
    -- CP-element group 771:  members (6) 
      -- CP-element group 771: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_sample_completed_
      -- CP-element group 771: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_update_start_
      -- CP-element group 771: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/$exit
      -- CP-element group 771: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/ack
      -- CP-element group 771: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/$entry
      -- CP-element group 771: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/req
      -- 
    ack_3508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 771_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1622_inst_ack_0, ack => concat_CP_34_elements(771)); -- 
    req_3512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(771), ack => WPIPE_Concat_output_pipe_1622_inst_req_1); -- 
    -- CP-element group 772:  transition  input  bypass 
    -- CP-element group 772: predecessors 
    -- CP-element group 772: 	771 
    -- CP-element group 772: successors 
    -- CP-element group 772: 	773 
    -- CP-element group 772:  members (3) 
      -- CP-element group 772: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_update_completed_
      -- CP-element group 772: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/$exit
      -- CP-element group 772: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/ack
      -- 
    ack_3513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 772_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1622_inst_ack_1, ack => concat_CP_34_elements(772)); -- 
    -- CP-element group 773:  join  transition  output  bypass 
    -- CP-element group 773: predecessors 
    -- CP-element group 773: 	763 
    -- CP-element group 773: 	772 
    -- CP-element group 773: successors 
    -- CP-element group 773: 	774 
    -- CP-element group 773:  members (3) 
      -- CP-element group 773: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_sample_start_
      -- CP-element group 773: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/$entry
      -- CP-element group 773: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/req
      -- 
    req_3521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(773), ack => WPIPE_Concat_output_pipe_1625_inst_req_0); -- 
    concat_cp_element_group_773: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_773"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(763) & concat_CP_34_elements(772);
      gj_concat_cp_element_group_773 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(773), clk => clk, reset => reset); --
    end block;
    -- CP-element group 774:  transition  input  output  bypass 
    -- CP-element group 774: predecessors 
    -- CP-element group 774: 	773 
    -- CP-element group 774: successors 
    -- CP-element group 774: 	775 
    -- CP-element group 774:  members (6) 
      -- CP-element group 774: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_sample_completed_
      -- CP-element group 774: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_update_start_
      -- CP-element group 774: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/$exit
      -- CP-element group 774: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/ack
      -- CP-element group 774: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/$entry
      -- CP-element group 774: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/req
      -- 
    ack_3522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 774_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1625_inst_ack_0, ack => concat_CP_34_elements(774)); -- 
    req_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(774), ack => WPIPE_Concat_output_pipe_1625_inst_req_1); -- 
    -- CP-element group 775:  transition  input  bypass 
    -- CP-element group 775: predecessors 
    -- CP-element group 775: 	774 
    -- CP-element group 775: successors 
    -- CP-element group 775: 	776 
    -- CP-element group 775:  members (3) 
      -- CP-element group 775: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_update_completed_
      -- CP-element group 775: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/$exit
      -- CP-element group 775: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/ack
      -- 
    ack_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 775_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1625_inst_ack_1, ack => concat_CP_34_elements(775)); -- 
    -- CP-element group 776:  join  transition  output  bypass 
    -- CP-element group 776: predecessors 
    -- CP-element group 776: 	761 
    -- CP-element group 776: 	775 
    -- CP-element group 776: successors 
    -- CP-element group 776: 	777 
    -- CP-element group 776:  members (3) 
      -- CP-element group 776: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_sample_start_
      -- CP-element group 776: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/$entry
      -- CP-element group 776: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/req
      -- 
    req_3535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(776), ack => WPIPE_Concat_output_pipe_1628_inst_req_0); -- 
    concat_cp_element_group_776: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_776"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(761) & concat_CP_34_elements(775);
      gj_concat_cp_element_group_776 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(776), clk => clk, reset => reset); --
    end block;
    -- CP-element group 777:  transition  input  output  bypass 
    -- CP-element group 777: predecessors 
    -- CP-element group 777: 	776 
    -- CP-element group 777: successors 
    -- CP-element group 777: 	778 
    -- CP-element group 777:  members (6) 
      -- CP-element group 777: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_sample_completed_
      -- CP-element group 777: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_update_start_
      -- CP-element group 777: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/$exit
      -- CP-element group 777: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/ack
      -- CP-element group 777: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/$entry
      -- CP-element group 777: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/req
      -- 
    ack_3536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 777_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1628_inst_ack_0, ack => concat_CP_34_elements(777)); -- 
    req_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(777), ack => WPIPE_Concat_output_pipe_1628_inst_req_1); -- 
    -- CP-element group 778:  transition  input  bypass 
    -- CP-element group 778: predecessors 
    -- CP-element group 778: 	777 
    -- CP-element group 778: successors 
    -- CP-element group 778: 	779 
    -- CP-element group 778:  members (3) 
      -- CP-element group 778: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_update_completed_
      -- CP-element group 778: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/$exit
      -- CP-element group 778: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/ack
      -- 
    ack_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 778_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1628_inst_ack_1, ack => concat_CP_34_elements(778)); -- 
    -- CP-element group 779:  join  transition  output  bypass 
    -- CP-element group 779: predecessors 
    -- CP-element group 779: 	759 
    -- CP-element group 779: 	778 
    -- CP-element group 779: successors 
    -- CP-element group 779: 	780 
    -- CP-element group 779:  members (3) 
      -- CP-element group 779: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_sample_start_
      -- CP-element group 779: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/$entry
      -- CP-element group 779: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/req
      -- 
    req_3549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(779), ack => WPIPE_Concat_output_pipe_1631_inst_req_0); -- 
    concat_cp_element_group_779: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_779"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(759) & concat_CP_34_elements(778);
      gj_concat_cp_element_group_779 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(779), clk => clk, reset => reset); --
    end block;
    -- CP-element group 780:  transition  input  output  bypass 
    -- CP-element group 780: predecessors 
    -- CP-element group 780: 	779 
    -- CP-element group 780: successors 
    -- CP-element group 780: 	781 
    -- CP-element group 780:  members (6) 
      -- CP-element group 780: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_sample_completed_
      -- CP-element group 780: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_update_start_
      -- CP-element group 780: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/$exit
      -- CP-element group 780: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/ack
      -- CP-element group 780: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/$entry
      -- CP-element group 780: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/req
      -- 
    ack_3550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 780_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1631_inst_ack_0, ack => concat_CP_34_elements(780)); -- 
    req_3554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(780), ack => WPIPE_Concat_output_pipe_1631_inst_req_1); -- 
    -- CP-element group 781:  transition  input  bypass 
    -- CP-element group 781: predecessors 
    -- CP-element group 781: 	780 
    -- CP-element group 781: successors 
    -- CP-element group 781: 	782 
    -- CP-element group 781:  members (3) 
      -- CP-element group 781: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_update_completed_
      -- CP-element group 781: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/$exit
      -- CP-element group 781: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/ack
      -- 
    ack_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 781_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1631_inst_ack_1, ack => concat_CP_34_elements(781)); -- 
    -- CP-element group 782:  join  transition  output  bypass 
    -- CP-element group 782: predecessors 
    -- CP-element group 782: 	757 
    -- CP-element group 782: 	781 
    -- CP-element group 782: successors 
    -- CP-element group 782: 	783 
    -- CP-element group 782:  members (3) 
      -- CP-element group 782: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_sample_start_
      -- CP-element group 782: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/$entry
      -- CP-element group 782: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/req
      -- 
    req_3563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(782), ack => WPIPE_Concat_output_pipe_1634_inst_req_0); -- 
    concat_cp_element_group_782: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_782"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(757) & concat_CP_34_elements(781);
      gj_concat_cp_element_group_782 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(782), clk => clk, reset => reset); --
    end block;
    -- CP-element group 783:  transition  input  output  bypass 
    -- CP-element group 783: predecessors 
    -- CP-element group 783: 	782 
    -- CP-element group 783: successors 
    -- CP-element group 783: 	784 
    -- CP-element group 783:  members (6) 
      -- CP-element group 783: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_sample_completed_
      -- CP-element group 783: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_update_start_
      -- CP-element group 783: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/$exit
      -- CP-element group 783: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/ack
      -- CP-element group 783: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/$entry
      -- CP-element group 783: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/req
      -- 
    ack_3564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 783_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1634_inst_ack_0, ack => concat_CP_34_elements(783)); -- 
    req_3568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(783), ack => WPIPE_Concat_output_pipe_1634_inst_req_1); -- 
    -- CP-element group 784:  transition  input  bypass 
    -- CP-element group 784: predecessors 
    -- CP-element group 784: 	783 
    -- CP-element group 784: successors 
    -- CP-element group 784: 	785 
    -- CP-element group 784:  members (3) 
      -- CP-element group 784: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_update_completed_
      -- CP-element group 784: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/$exit
      -- CP-element group 784: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/ack
      -- 
    ack_3569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 784_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1634_inst_ack_1, ack => concat_CP_34_elements(784)); -- 
    -- CP-element group 785:  join  transition  output  bypass 
    -- CP-element group 785: predecessors 
    -- CP-element group 785: 	755 
    -- CP-element group 785: 	784 
    -- CP-element group 785: successors 
    -- CP-element group 785: 	786 
    -- CP-element group 785:  members (3) 
      -- CP-element group 785: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_sample_start_
      -- CP-element group 785: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/$entry
      -- CP-element group 785: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/req
      -- 
    req_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(785), ack => WPIPE_Concat_output_pipe_1637_inst_req_0); -- 
    concat_cp_element_group_785: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_785"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(755) & concat_CP_34_elements(784);
      gj_concat_cp_element_group_785 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(785), clk => clk, reset => reset); --
    end block;
    -- CP-element group 786:  transition  input  output  bypass 
    -- CP-element group 786: predecessors 
    -- CP-element group 786: 	785 
    -- CP-element group 786: successors 
    -- CP-element group 786: 	787 
    -- CP-element group 786:  members (6) 
      -- CP-element group 786: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_sample_completed_
      -- CP-element group 786: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_update_start_
      -- CP-element group 786: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/$exit
      -- CP-element group 786: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/ack
      -- CP-element group 786: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/$entry
      -- CP-element group 786: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/req
      -- 
    ack_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 786_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1637_inst_ack_0, ack => concat_CP_34_elements(786)); -- 
    req_3582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(786), ack => WPIPE_Concat_output_pipe_1637_inst_req_1); -- 
    -- CP-element group 787:  transition  input  bypass 
    -- CP-element group 787: predecessors 
    -- CP-element group 787: 	786 
    -- CP-element group 787: successors 
    -- CP-element group 787: 	788 
    -- CP-element group 787:  members (3) 
      -- CP-element group 787: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_update_completed_
      -- CP-element group 787: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/$exit
      -- CP-element group 787: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/ack
      -- 
    ack_3583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 787_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1637_inst_ack_1, ack => concat_CP_34_elements(787)); -- 
    -- CP-element group 788:  join  transition  output  bypass 
    -- CP-element group 788: predecessors 
    -- CP-element group 788: 	753 
    -- CP-element group 788: 	787 
    -- CP-element group 788: successors 
    -- CP-element group 788: 	789 
    -- CP-element group 788:  members (3) 
      -- CP-element group 788: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_sample_start_
      -- CP-element group 788: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/$entry
      -- CP-element group 788: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/req
      -- 
    req_3591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(788), ack => WPIPE_Concat_output_pipe_1640_inst_req_0); -- 
    concat_cp_element_group_788: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_788"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(753) & concat_CP_34_elements(787);
      gj_concat_cp_element_group_788 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(788), clk => clk, reset => reset); --
    end block;
    -- CP-element group 789:  transition  input  output  bypass 
    -- CP-element group 789: predecessors 
    -- CP-element group 789: 	788 
    -- CP-element group 789: successors 
    -- CP-element group 789: 	790 
    -- CP-element group 789:  members (6) 
      -- CP-element group 789: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_sample_completed_
      -- CP-element group 789: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_update_start_
      -- CP-element group 789: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/$exit
      -- CP-element group 789: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/ack
      -- CP-element group 789: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/$entry
      -- CP-element group 789: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/req
      -- 
    ack_3592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 789_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1640_inst_ack_0, ack => concat_CP_34_elements(789)); -- 
    req_3596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(789), ack => WPIPE_Concat_output_pipe_1640_inst_req_1); -- 
    -- CP-element group 790:  transition  input  bypass 
    -- CP-element group 790: predecessors 
    -- CP-element group 790: 	789 
    -- CP-element group 790: successors 
    -- CP-element group 790: 	791 
    -- CP-element group 790:  members (3) 
      -- CP-element group 790: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_update_completed_
      -- CP-element group 790: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/$exit
      -- CP-element group 790: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/ack
      -- 
    ack_3597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 790_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1640_inst_ack_1, ack => concat_CP_34_elements(790)); -- 
    -- CP-element group 791:  branch  join  transition  place  output  bypass 
    -- CP-element group 791: predecessors 
    -- CP-element group 791: 	746 
    -- CP-element group 791: 	790 
    -- CP-element group 791: successors 
    -- CP-element group 791: 	792 
    -- CP-element group 791: 	793 
    -- CP-element group 791:  members (10) 
      -- CP-element group 791: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653__exit__
      -- CP-element group 791: 	 branch_block_stmt_23/if_stmt_1654__entry__
      -- CP-element group 791: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/$exit
      -- CP-element group 791: 	 branch_block_stmt_23/if_stmt_1654_dead_link/$entry
      -- CP-element group 791: 	 branch_block_stmt_23/if_stmt_1654_eval_test/$entry
      -- CP-element group 791: 	 branch_block_stmt_23/if_stmt_1654_eval_test/$exit
      -- CP-element group 791: 	 branch_block_stmt_23/if_stmt_1654_eval_test/branch_req
      -- CP-element group 791: 	 branch_block_stmt_23/R_exitcond1_1655_place
      -- CP-element group 791: 	 branch_block_stmt_23/if_stmt_1654_if_link/$entry
      -- CP-element group 791: 	 branch_block_stmt_23/if_stmt_1654_else_link/$entry
      -- 
    branch_req_3605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(791), ack => if_stmt_1654_branch_req_0); -- 
    concat_cp_element_group_791: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_791"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(746) & concat_CP_34_elements(790);
      gj_concat_cp_element_group_791 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(791), clk => clk, reset => reset); --
    end block;
    -- CP-element group 792:  merge  transition  place  input  bypass 
    -- CP-element group 792: predecessors 
    -- CP-element group 792: 	791 
    -- CP-element group 792: successors 
    -- CP-element group 792: 	802 
    -- CP-element group 792:  members (13) 
      -- CP-element group 792: 	 branch_block_stmt_23/merge_stmt_1660__exit__
      -- CP-element group 792: 	 branch_block_stmt_23/forx_xend453x_xloopexit_forx_xend453
      -- CP-element group 792: 	 branch_block_stmt_23/if_stmt_1654_if_link/$exit
      -- CP-element group 792: 	 branch_block_stmt_23/if_stmt_1654_if_link/if_choice_transition
      -- CP-element group 792: 	 branch_block_stmt_23/forx_xbody380_forx_xend453x_xloopexit
      -- CP-element group 792: 	 branch_block_stmt_23/forx_xbody380_forx_xend453x_xloopexit_PhiReq/$entry
      -- CP-element group 792: 	 branch_block_stmt_23/forx_xbody380_forx_xend453x_xloopexit_PhiReq/$exit
      -- CP-element group 792: 	 branch_block_stmt_23/merge_stmt_1660_PhiReqMerge
      -- CP-element group 792: 	 branch_block_stmt_23/merge_stmt_1660_PhiAck/$entry
      -- CP-element group 792: 	 branch_block_stmt_23/merge_stmt_1660_PhiAck/$exit
      -- CP-element group 792: 	 branch_block_stmt_23/merge_stmt_1660_PhiAck/dummy
      -- CP-element group 792: 	 branch_block_stmt_23/forx_xend453x_xloopexit_forx_xend453_PhiReq/$entry
      -- CP-element group 792: 	 branch_block_stmt_23/forx_xend453x_xloopexit_forx_xend453_PhiReq/$exit
      -- 
    if_choice_transition_3610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 792_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1654_branch_ack_1, ack => concat_CP_34_elements(792)); -- 
    -- CP-element group 793:  fork  transition  place  input  output  bypass 
    -- CP-element group 793: predecessors 
    -- CP-element group 793: 	791 
    -- CP-element group 793: successors 
    -- CP-element group 793: 	797 
    -- CP-element group 793: 	798 
    -- CP-element group 793:  members (12) 
      -- CP-element group 793: 	 branch_block_stmt_23/if_stmt_1654_else_link/$exit
      -- CP-element group 793: 	 branch_block_stmt_23/if_stmt_1654_else_link/else_choice_transition
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/$entry
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/$entry
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$entry
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/$entry
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/$entry
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/$entry
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/rr
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/$entry
      -- CP-element group 793: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 793_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1654_branch_ack_0, ack => concat_CP_34_elements(793)); -- 
    rr_3761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(793), ack => type_cast_1532_inst_req_0); -- 
    cr_3766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(793), ack => type_cast_1532_inst_req_1); -- 
    -- CP-element group 794:  merge  branch  transition  place  output  bypass 
    -- CP-element group 794: predecessors 
    -- CP-element group 794: 	78 
    -- CP-element group 794: 	192 
    -- CP-element group 794: successors 
    -- CP-element group 794: 	79 
    -- CP-element group 794: 	80 
    -- CP-element group 794:  members (17) 
      -- CP-element group 794: 	 branch_block_stmt_23/merge_stmt_306__exit__
      -- CP-element group 794: 	 branch_block_stmt_23/assign_stmt_312__entry__
      -- CP-element group 794: 	 branch_block_stmt_23/assign_stmt_312__exit__
      -- CP-element group 794: 	 branch_block_stmt_23/if_stmt_313__entry__
      -- CP-element group 794: 	 branch_block_stmt_23/assign_stmt_312/$entry
      -- CP-element group 794: 	 branch_block_stmt_23/assign_stmt_312/$exit
      -- CP-element group 794: 	 branch_block_stmt_23/if_stmt_313_dead_link/$entry
      -- CP-element group 794: 	 branch_block_stmt_23/if_stmt_313_eval_test/$entry
      -- CP-element group 794: 	 branch_block_stmt_23/if_stmt_313_eval_test/$exit
      -- CP-element group 794: 	 branch_block_stmt_23/if_stmt_313_eval_test/branch_req
      -- CP-element group 794: 	 branch_block_stmt_23/R_cmp167463_314_place
      -- CP-element group 794: 	 branch_block_stmt_23/if_stmt_313_if_link/$entry
      -- CP-element group 794: 	 branch_block_stmt_23/if_stmt_313_else_link/$entry
      -- CP-element group 794: 	 branch_block_stmt_23/merge_stmt_306_PhiReqMerge
      -- CP-element group 794: 	 branch_block_stmt_23/merge_stmt_306_PhiAck/$entry
      -- CP-element group 794: 	 branch_block_stmt_23/merge_stmt_306_PhiAck/$exit
      -- CP-element group 794: 	 branch_block_stmt_23/merge_stmt_306_PhiAck/dummy
      -- 
    branch_req_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(794), ack => if_stmt_313_branch_req_0); -- 
    concat_CP_34_elements(794) <= OrReduce(concat_CP_34_elements(78) & concat_CP_34_elements(192));
    -- CP-element group 795:  merge  fork  transition  place  output  bypass 
    -- CP-element group 795: predecessors 
    -- CP-element group 795: 	80 
    -- CP-element group 795: 	305 
    -- CP-element group 795: successors 
    -- CP-element group 795: 	307 
    -- CP-element group 795: 	308 
    -- CP-element group 795:  members (13) 
      -- CP-element group 795: 	 branch_block_stmt_23/merge_stmt_765__exit__
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768__entry__
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768/$entry
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_sample_start_
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_update_start_
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/$entry
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/crr
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/$entry
      -- CP-element group 795: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/ccr
      -- CP-element group 795: 	 branch_block_stmt_23/merge_stmt_765_PhiReqMerge
      -- CP-element group 795: 	 branch_block_stmt_23/merge_stmt_765_PhiAck/$entry
      -- CP-element group 795: 	 branch_block_stmt_23/merge_stmt_765_PhiAck/$exit
      -- CP-element group 795: 	 branch_block_stmt_23/merge_stmt_765_PhiAck/dummy
      -- 
    crr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(795), ack => call_stmt_768_call_req_0); -- 
    ccr_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(795), ack => call_stmt_768_call_req_1); -- 
    concat_CP_34_elements(795) <= OrReduce(concat_CP_34_elements(80) & concat_CP_34_elements(305));
    -- CP-element group 796:  transition  output  delay-element  bypass 
    -- CP-element group 796: predecessors 
    -- CP-element group 796: 	745 
    -- CP-element group 796: successors 
    -- CP-element group 796: 	800 
    -- CP-element group 796:  members (5) 
      -- CP-element group 796: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/$exit
      -- CP-element group 796: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/phi_stmt_1526/$exit
      -- CP-element group 796: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$exit
      -- CP-element group 796: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1530_konst_delay_trans
      -- CP-element group 796: 	 branch_block_stmt_23/bbx_xnph_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_req
      -- 
    phi_stmt_1526_req_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1526_req_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(796), ack => phi_stmt_1526_req_0); -- 
    -- Element group concat_CP_34_elements(796) is a control-delay.
    cp_element_796_delay: control_delay_element  generic map(name => " 796_delay", delay_value => 1)  port map(req => concat_CP_34_elements(745), ack => concat_CP_34_elements(796), clk => clk, reset =>reset);
    -- CP-element group 797:  transition  input  bypass 
    -- CP-element group 797: predecessors 
    -- CP-element group 797: 	793 
    -- CP-element group 797: successors 
    -- CP-element group 797: 	799 
    -- CP-element group 797:  members (2) 
      -- CP-element group 797: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/$exit
      -- CP-element group 797: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/ra
      -- 
    ra_3762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 797_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1532_inst_ack_0, ack => concat_CP_34_elements(797)); -- 
    -- CP-element group 798:  transition  input  bypass 
    -- CP-element group 798: predecessors 
    -- CP-element group 798: 	793 
    -- CP-element group 798: successors 
    -- CP-element group 798: 	799 
    -- CP-element group 798:  members (2) 
      -- CP-element group 798: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/$exit
      -- CP-element group 798: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/ca
      -- 
    ca_3767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 798_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1532_inst_ack_1, ack => concat_CP_34_elements(798)); -- 
    -- CP-element group 799:  join  transition  output  bypass 
    -- CP-element group 799: predecessors 
    -- CP-element group 799: 	797 
    -- CP-element group 799: 	798 
    -- CP-element group 799: successors 
    -- CP-element group 799: 	800 
    -- CP-element group 799:  members (6) 
      -- CP-element group 799: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/$exit
      -- CP-element group 799: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/$exit
      -- CP-element group 799: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$exit
      -- CP-element group 799: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/$exit
      -- CP-element group 799: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/$exit
      -- CP-element group 799: 	 branch_block_stmt_23/forx_xbody380_forx_xbody380_PhiReq/phi_stmt_1526/phi_stmt_1526_req
      -- 
    phi_stmt_1526_req_3768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1526_req_3768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(799), ack => phi_stmt_1526_req_1); -- 
    concat_cp_element_group_799: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_799"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(797) & concat_CP_34_elements(798);
      gj_concat_cp_element_group_799 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(799), clk => clk, reset => reset); --
    end block;
    -- CP-element group 800:  merge  transition  place  bypass 
    -- CP-element group 800: predecessors 
    -- CP-element group 800: 	796 
    -- CP-element group 800: 	799 
    -- CP-element group 800: successors 
    -- CP-element group 800: 	801 
    -- CP-element group 800:  members (2) 
      -- CP-element group 800: 	 branch_block_stmt_23/merge_stmt_1525_PhiReqMerge
      -- CP-element group 800: 	 branch_block_stmt_23/merge_stmt_1525_PhiAck/$entry
      -- 
    concat_CP_34_elements(800) <= OrReduce(concat_CP_34_elements(796) & concat_CP_34_elements(799));
    -- CP-element group 801:  fork  transition  place  input  output  bypass 
    -- CP-element group 801: predecessors 
    -- CP-element group 801: 	800 
    -- CP-element group 801: successors 
    -- CP-element group 801: 	746 
    -- CP-element group 801: 	747 
    -- CP-element group 801: 	749 
    -- CP-element group 801: 	751 
    -- CP-element group 801: 	753 
    -- CP-element group 801: 	755 
    -- CP-element group 801: 	757 
    -- CP-element group 801: 	759 
    -- CP-element group 801: 	761 
    -- CP-element group 801: 	763 
    -- CP-element group 801: 	765 
    -- CP-element group 801: 	767 
    -- CP-element group 801:  members (53) 
      -- CP-element group 801: 	 branch_block_stmt_23/merge_stmt_1525__exit__
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653__entry__
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/req
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/req
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resized_1
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scaled_1
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_computed_1
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/$exit
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/index_resize_req
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/index_resize_ack
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/$exit
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/scale_rename_req
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/scale_rename_ack
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_update_start
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/req
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_update_start_
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/cr
      -- CP-element group 801: 	 branch_block_stmt_23/merge_stmt_1525_PhiAck/$exit
      -- CP-element group 801: 	 branch_block_stmt_23/merge_stmt_1525_PhiAck/phi_stmt_1526_ack
      -- 
    phi_stmt_1526_ack_3773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 801_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1526_ack_0, ack => concat_CP_34_elements(801)); -- 
    req_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => array_obj_ref_1538_index_offset_req_0); -- 
    cr_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1597_inst_req_1); -- 
    req_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => array_obj_ref_1538_index_offset_req_1); -- 
    cr_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1587_inst_req_1); -- 
    cr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1567_inst_req_1); -- 
    cr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1547_inst_req_1); -- 
    cr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => ptr_deref_1543_load_0_req_1); -- 
    cr_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1557_inst_req_1); -- 
    req_3322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => addr_of_1539_final_reg_req_1); -- 
    cr_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1577_inst_req_1); -- 
    cr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1607_inst_req_1); -- 
    cr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(801), ack => type_cast_1617_inst_req_1); -- 
    -- CP-element group 802:  merge  transition  place  bypass 
    -- CP-element group 802: predecessors 
    -- CP-element group 802: 	743 
    -- CP-element group 802: 	792 
    -- CP-element group 802: successors 
    -- CP-element group 802:  members (16) 
      -- CP-element group 802: 	 $exit
      -- CP-element group 802: 	 branch_block_stmt_23/$exit
      -- CP-element group 802: 	 branch_block_stmt_23/branch_block_stmt_23__exit__
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1662__exit__
      -- CP-element group 802: 	 branch_block_stmt_23/return__
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1664__exit__
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1662_PhiReqMerge
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1662_PhiAck/$entry
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1662_PhiAck/$exit
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1662_PhiAck/dummy
      -- CP-element group 802: 	 branch_block_stmt_23/return___PhiReq/$entry
      -- CP-element group 802: 	 branch_block_stmt_23/return___PhiReq/$exit
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1664_PhiReqMerge
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1664_PhiAck/$entry
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1664_PhiAck/$exit
      -- CP-element group 802: 	 branch_block_stmt_23/merge_stmt_1664_PhiAck/dummy
      -- 
    concat_CP_34_elements(802) <= OrReduce(concat_CP_34_elements(743) & concat_CP_34_elements(792));
    concat_do_while_stmt_368_terminator_1072: loop_terminator -- 
      generic map (name => " concat_do_while_stmt_368_terminator_1072", max_iterations_in_flight =>15) 
      port map(loop_body_exit => concat_CP_34_elements(87),loop_continue => concat_CP_34_elements(190),loop_terminate => concat_CP_34_elements(189),loop_back => concat_CP_34_elements(85),loop_exit => concat_CP_34_elements(84),clk => clk, reset => reset); -- 
    phi_stmt_370_phi_seq_742_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(97);
      concat_CP_34_elements(102)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(106);
      concat_CP_34_elements(103)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(107);
      concat_CP_34_elements(98) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(99);
      concat_CP_34_elements(108)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(108);
      concat_CP_34_elements(109)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(110);
      concat_CP_34_elements(100) <= phi_mux_reqs(1);
      phi_stmt_370_phi_seq_742 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_370_phi_seq_742") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(92), 
          phi_sample_ack => concat_CP_34_elements(95), 
          phi_update_req => concat_CP_34_elements(94), 
          phi_update_ack => concat_CP_34_elements(96), 
          phi_mux_ack => concat_CP_34_elements(101), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_694_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= concat_CP_34_elements(88);
        preds(1)  <= concat_CP_34_elements(89);
        entry_tmerge_694 : transition_merge -- 
          generic map(name => " entry_tmerge_694")
          port map (preds => preds, symbol_out => concat_CP_34_elements(90));
          -- 
    end block;
    concat_do_while_stmt_590_terminator_1501: loop_terminator -- 
      generic map (name => " concat_do_while_stmt_590_terminator_1501", max_iterations_in_flight =>15) 
      port map(loop_body_exit => concat_CP_34_elements(200),loop_continue => concat_CP_34_elements(303),loop_terminate => concat_CP_34_elements(302),loop_back => concat_CP_34_elements(198),loop_exit => concat_CP_34_elements(197),clk => clk, reset => reset); -- 
    phi_stmt_592_phi_seq_1171_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(210);
      concat_CP_34_elements(215)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(219);
      concat_CP_34_elements(216)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(220);
      concat_CP_34_elements(211) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(212);
      concat_CP_34_elements(221)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(221);
      concat_CP_34_elements(222)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(223);
      concat_CP_34_elements(213) <= phi_mux_reqs(1);
      phi_stmt_592_phi_seq_1171 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_592_phi_seq_1171") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(205), 
          phi_sample_ack => concat_CP_34_elements(208), 
          phi_update_req => concat_CP_34_elements(207), 
          phi_update_ack => concat_CP_34_elements(209), 
          phi_mux_ack => concat_CP_34_elements(214), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1123_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= concat_CP_34_elements(201);
        preds(1)  <= concat_CP_34_elements(202);
        entry_tmerge_1123 : transition_merge -- 
          generic map(name => " entry_tmerge_1123")
          port map (preds => preds, symbol_out => concat_CP_34_elements(203));
          -- 
    end block;
    concat_do_while_stmt_817_terminator_2945: loop_terminator -- 
      generic map (name => " concat_do_while_stmt_817_terminator_2945", max_iterations_in_flight =>15) 
      port map(loop_body_exit => concat_CP_34_elements(313),loop_continue => concat_CP_34_elements(693),loop_terminate => concat_CP_34_elements(692),loop_back => concat_CP_34_elements(311),loop_exit => concat_CP_34_elements(310),clk => clk, reset => reset); -- 
    phi_stmt_819_phi_seq_1603_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(328);
      concat_CP_34_elements(333)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(337);
      concat_CP_34_elements(334)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(338);
      concat_CP_34_elements(329) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(330);
      concat_CP_34_elements(339)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(339);
      concat_CP_34_elements(340)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(341);
      concat_CP_34_elements(331) <= phi_mux_reqs(1);
      phi_stmt_819_phi_seq_1603 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_819_phi_seq_1603") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(324), 
          phi_sample_ack => concat_CP_34_elements(325), 
          phi_update_req => concat_CP_34_elements(326), 
          phi_update_ack => concat_CP_34_elements(327), 
          phi_mux_ack => concat_CP_34_elements(332), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_824_phi_seq_1647_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(347);
      concat_CP_34_elements(352)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(356);
      concat_CP_34_elements(353)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(357);
      concat_CP_34_elements(348) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(349);
      concat_CP_34_elements(358)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(358);
      concat_CP_34_elements(359)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(360);
      concat_CP_34_elements(350) <= phi_mux_reqs(1);
      phi_stmt_824_phi_seq_1647 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_824_phi_seq_1647") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(318), 
          phi_sample_ack => concat_CP_34_elements(345), 
          phi_update_req => concat_CP_34_elements(320), 
          phi_update_ack => concat_CP_34_elements(346), 
          phi_mux_ack => concat_CP_34_elements(351), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_829_phi_seq_1691_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(368);
      concat_CP_34_elements(373)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(377);
      concat_CP_34_elements(374)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(378);
      concat_CP_34_elements(369) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(370);
      concat_CP_34_elements(379)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(379);
      concat_CP_34_elements(380)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(381);
      concat_CP_34_elements(371) <= phi_mux_reqs(1);
      phi_stmt_829_phi_seq_1691 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_829_phi_seq_1691") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(364), 
          phi_sample_ack => concat_CP_34_elements(365), 
          phi_update_req => concat_CP_34_elements(366), 
          phi_update_ack => concat_CP_34_elements(367), 
          phi_mux_ack => concat_CP_34_elements(372), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_834_phi_seq_1735_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(389);
      concat_CP_34_elements(394)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(398);
      concat_CP_34_elements(395)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(399);
      concat_CP_34_elements(390) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(391);
      concat_CP_34_elements(400)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(400);
      concat_CP_34_elements(401)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(402);
      concat_CP_34_elements(392) <= phi_mux_reqs(1);
      phi_stmt_834_phi_seq_1735 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_834_phi_seq_1735") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(385), 
          phi_sample_ack => concat_CP_34_elements(386), 
          phi_update_req => concat_CP_34_elements(387), 
          phi_update_ack => concat_CP_34_elements(388), 
          phi_mux_ack => concat_CP_34_elements(393), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_839_phi_seq_1779_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(410);
      concat_CP_34_elements(415)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(419);
      concat_CP_34_elements(416)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(420);
      concat_CP_34_elements(411) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(412);
      concat_CP_34_elements(421)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(421);
      concat_CP_34_elements(422)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(423);
      concat_CP_34_elements(413) <= phi_mux_reqs(1);
      phi_stmt_839_phi_seq_1779 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_839_phi_seq_1779") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(406), 
          phi_sample_ack => concat_CP_34_elements(407), 
          phi_update_req => concat_CP_34_elements(408), 
          phi_update_ack => concat_CP_34_elements(409), 
          phi_mux_ack => concat_CP_34_elements(414), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1555_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= concat_CP_34_elements(314);
        preds(1)  <= concat_CP_34_elements(315);
        entry_tmerge_1555 : transition_merge -- 
          generic map(name => " entry_tmerge_1555")
          port map (preds => preds, symbol_out => concat_CP_34_elements(316));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_1152_1152_delayed_2_0_1254 : std_logic_vector(15 downto 0);
    signal MUX_1166_wire : std_logic_vector(15 downto 0);
    signal MUX_1168_1168_delayed_2_0_1282 : std_logic_vector(15 downto 0);
    signal MUX_1181_wire : std_logic_vector(15 downto 0);
    signal MUX_1185_1185_delayed_2_0_1306 : std_logic_vector(15 downto 0);
    signal MUX_1196_wire : std_logic_vector(15 downto 0);
    signal MUX_1202_1202_delayed_2_0_1332 : std_logic_vector(15 downto 0);
    signal MUX_1261_wire : std_logic_vector(15 downto 0);
    signal MUX_1289_wire : std_logic_vector(15 downto 0);
    signal MUX_1315_wire : std_logic_vector(15 downto 0);
    signal MUX_1341_wire : std_logic_vector(15 downto 0);
    signal MUX_963_wire : std_logic_vector(15 downto 0);
    signal MUX_978_wire : std_logic_vector(15 downto 0);
    signal MUX_993_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1024_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1061_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1227_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1358_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_536_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_758_wire : std_logic_vector(0 downto 0);
    signal R_idxprom240_875_resized : std_logic_vector(13 downto 0);
    signal R_idxprom240_875_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom244_898_resized : std_logic_vector(13 downto 0);
    signal R_idxprom244_898_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom268_1078_resized : std_logic_vector(13 downto 0);
    signal R_idxprom268_1078_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom272_1101_resized : std_logic_vector(13 downto 0);
    signal R_idxprom272_1101_scaled : std_logic_vector(13 downto 0);
    signal R_indvar476_601_resized : std_logic_vector(13 downto 0);
    signal R_indvar476_601_scaled : std_logic_vector(13 downto 0);
    signal R_indvar488_379_resized : std_logic_vector(13 downto 0);
    signal R_indvar488_379_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1537_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1537_scaled : std_logic_vector(13 downto 0);
    signal add123_407 : std_logic_vector(63 downto 0);
    signal add129_425 : std_logic_vector(63 downto 0);
    signal add12_74 : std_logic_vector(31 downto 0);
    signal add135_443 : std_logic_vector(63 downto 0);
    signal add141_461 : std_logic_vector(63 downto 0);
    signal add147_479 : std_logic_vector(63 downto 0);
    signal add153_497 : std_logic_vector(63 downto 0);
    signal add159_515 : std_logic_vector(63 downto 0);
    signal add179_629 : std_logic_vector(63 downto 0);
    signal add185_647 : std_logic_vector(63 downto 0);
    signal add191_665 : std_logic_vector(63 downto 0);
    signal add197_683 : std_logic_vector(63 downto 0);
    signal add203_701 : std_logic_vector(63 downto 0);
    signal add209_719 : std_logic_vector(63 downto 0);
    signal add215_737 : std_logic_vector(63 downto 0);
    signal add21_99 : std_logic_vector(31 downto 0);
    signal add30_124 : std_logic_vector(31 downto 0);
    signal add39_149 : std_logic_vector(31 downto 0);
    signal add48_174 : std_logic_vector(31 downto 0);
    signal add57_199 : std_logic_vector(31 downto 0);
    signal add66_224 : std_logic_vector(31 downto 0);
    signal add75_249 : std_logic_vector(31 downto 0);
    signal add_49 : std_logic_vector(31 downto 0);
    signal add_inp1x_x0_980 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_824 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_866_delayed_1_0_866 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_907_delayed_1_0_925 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_at_entry_796 : std_logic_vector(15 downto 0);
    signal add_inp2x_x0504_1263 : std_logic_vector(15 downto 0);
    signal add_inp2x_x0x_xph_1183 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_1015_delayed_3_0_1069 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_1056_delayed_3_0_1128 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_829 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_at_entry_801 : std_logic_vector(15 downto 0);
    signal add_outx_x0_1032_delayed_2_0_1092 : std_logic_vector(15 downto 0);
    signal add_outx_x0_1063_delayed_2_0_1138 : std_logic_vector(15 downto 0);
    signal add_outx_x0_965 : std_logic_vector(15 downto 0);
    signal add_outx_x1_819 : std_logic_vector(15 downto 0);
    signal add_outx_x1_883_delayed_1_0_889 : std_logic_vector(15 downto 0);
    signal add_outx_x1_914_delayed_1_0_935 : std_logic_vector(15 downto 0);
    signal add_outx_x1_at_entry_790 : std_logic_vector(15 downto 0);
    signal add_outx_x2502_1291 : std_logic_vector(15 downto 0);
    signal add_outx_x2x_xph_1168 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1079_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_380_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_380_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_380_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_380_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_380_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_380_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_602_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_602_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_602_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_602_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_602_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_602_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_root_address : std_logic_vector(13 downto 0);
    signal arrayidx219_604 : std_logic_vector(31 downto 0);
    signal arrayidx241_878 : std_logic_vector(31 downto 0);
    signal arrayidx245_894_delayed_6_0_907 : std_logic_vector(31 downto 0);
    signal arrayidx245_901 : std_logic_vector(31 downto 0);
    signal arrayidx269_1081 : std_logic_vector(31 downto 0);
    signal arrayidx273_1043_delayed_6_0_1110 : std_logic_vector(31 downto 0);
    signal arrayidx273_1104 : std_logic_vector(31 downto 0);
    signal arrayidx385_1540 : std_logic_vector(31 downto 0);
    signal arrayidx_382 : std_logic_vector(31 downto 0);
    signal call10_65 : std_logic_vector(7 downto 0);
    signal call116_385 : std_logic_vector(7 downto 0);
    signal call120_398 : std_logic_vector(7 downto 0);
    signal call126_416 : std_logic_vector(7 downto 0);
    signal call132_434 : std_logic_vector(7 downto 0);
    signal call138_452 : std_logic_vector(7 downto 0);
    signal call144_470 : std_logic_vector(7 downto 0);
    signal call14_77 : std_logic_vector(7 downto 0);
    signal call150_488 : std_logic_vector(7 downto 0);
    signal call156_506 : std_logic_vector(7 downto 0);
    signal call172_607 : std_logic_vector(7 downto 0);
    signal call176_620 : std_logic_vector(7 downto 0);
    signal call182_638 : std_logic_vector(7 downto 0);
    signal call188_656 : std_logic_vector(7 downto 0);
    signal call194_674 : std_logic_vector(7 downto 0);
    signal call19_90 : std_logic_vector(7 downto 0);
    signal call200_692 : std_logic_vector(7 downto 0);
    signal call206_710 : std_logic_vector(7 downto 0);
    signal call212_728 : std_logic_vector(7 downto 0);
    signal call225_768 : std_logic_vector(63 downto 0);
    signal call23_102 : std_logic_vector(7 downto 0);
    signal call28_115 : std_logic_vector(7 downto 0);
    signal call2_40 : std_logic_vector(7 downto 0);
    signal call307_1372 : std_logic_vector(63 downto 0);
    signal call32_127 : std_logic_vector(7 downto 0);
    signal call37_140 : std_logic_vector(7 downto 0);
    signal call41_152 : std_logic_vector(7 downto 0);
    signal call46_165 : std_logic_vector(7 downto 0);
    signal call50_177 : std_logic_vector(7 downto 0);
    signal call55_190 : std_logic_vector(7 downto 0);
    signal call59_202 : std_logic_vector(7 downto 0);
    signal call5_52 : std_logic_vector(7 downto 0);
    signal call64_215 : std_logic_vector(7 downto 0);
    signal call68_227 : std_logic_vector(7 downto 0);
    signal call73_240 : std_logic_vector(7 downto 0);
    signal call_26 : std_logic_vector(7 downto 0);
    signal cmp167463_312 : std_logic_vector(0 downto 0);
    signal cmp237_853 : std_logic_vector(0 downto 0);
    signal cmp257_1009 : std_logic_vector(0 downto 0);
    signal cmp264_1046 : std_logic_vector(0 downto 0);
    signal cmp294_1212 : std_logic_vector(0 downto 0);
    signal cmp302_1352 : std_logic_vector(0 downto 0);
    signal cmp378460_1487 : std_logic_vector(0 downto 0);
    signal cmp467_297 : std_logic_vector(0 downto 0);
    signal conv102_275 : std_logic_vector(31 downto 0);
    signal conv108_286 : std_logic_vector(31 downto 0);
    signal conv117_389 : std_logic_vector(63 downto 0);
    signal conv11_69 : std_logic_vector(31 downto 0);
    signal conv122_402 : std_logic_vector(63 downto 0);
    signal conv128_420 : std_logic_vector(63 downto 0);
    signal conv134_438 : std_logic_vector(63 downto 0);
    signal conv140_456 : std_logic_vector(63 downto 0);
    signal conv146_474 : std_logic_vector(63 downto 0);
    signal conv152_492 : std_logic_vector(63 downto 0);
    signal conv158_510 : std_logic_vector(63 downto 0);
    signal conv173_611 : std_logic_vector(63 downto 0);
    signal conv178_624 : std_logic_vector(63 downto 0);
    signal conv17_81 : std_logic_vector(31 downto 0);
    signal conv184_642 : std_logic_vector(63 downto 0);
    signal conv190_660 : std_logic_vector(63 downto 0);
    signal conv196_678 : std_logic_vector(63 downto 0);
    signal conv1_31 : std_logic_vector(31 downto 0);
    signal conv202_696 : std_logic_vector(63 downto 0);
    signal conv208_714 : std_logic_vector(63 downto 0);
    signal conv20_94 : std_logic_vector(31 downto 0);
    signal conv214_732 : std_logic_vector(63 downto 0);
    signal conv226_1369 : std_logic_vector(63 downto 0);
    signal conv233_848 : std_logic_vector(31 downto 0);
    signal conv253_1000 : std_logic_vector(31 downto 0);
    signal conv260_1037 : std_logic_vector(31 downto 0);
    signal conv26_106 : std_logic_vector(31 downto 0);
    signal conv290_1203 : std_logic_vector(31 downto 0);
    signal conv299_1347 : std_logic_vector(31 downto 0);
    signal conv29_119 : std_logic_vector(31 downto 0);
    signal conv308_1377 : std_logic_vector(63 downto 0);
    signal conv314_1386 : std_logic_vector(7 downto 0);
    signal conv320_1396 : std_logic_vector(7 downto 0);
    signal conv326_1406 : std_logic_vector(7 downto 0);
    signal conv332_1416 : std_logic_vector(7 downto 0);
    signal conv338_1426 : std_logic_vector(7 downto 0);
    signal conv344_1436 : std_logic_vector(7 downto 0);
    signal conv350_1446 : std_logic_vector(7 downto 0);
    signal conv356_1456 : std_logic_vector(7 downto 0);
    signal conv35_131 : std_logic_vector(31 downto 0);
    signal conv38_144 : std_logic_vector(31 downto 0);
    signal conv390_1548 : std_logic_vector(7 downto 0);
    signal conv396_1558 : std_logic_vector(7 downto 0);
    signal conv3_44 : std_logic_vector(31 downto 0);
    signal conv402_1568 : std_logic_vector(7 downto 0);
    signal conv408_1578 : std_logic_vector(7 downto 0);
    signal conv414_1588 : std_logic_vector(7 downto 0);
    signal conv420_1598 : std_logic_vector(7 downto 0);
    signal conv426_1608 : std_logic_vector(7 downto 0);
    signal conv432_1618 : std_logic_vector(7 downto 0);
    signal conv44_156 : std_logic_vector(31 downto 0);
    signal conv47_169 : std_logic_vector(31 downto 0);
    signal conv53_181 : std_logic_vector(31 downto 0);
    signal conv56_194 : std_logic_vector(31 downto 0);
    signal conv62_206 : std_logic_vector(31 downto 0);
    signal conv65_219 : std_logic_vector(31 downto 0);
    signal conv71_231 : std_logic_vector(31 downto 0);
    signal conv74_244 : std_logic_vector(31 downto 0);
    signal conv8_56 : std_logic_vector(31 downto 0);
    signal count_inp1x_x0_995 : std_logic_vector(15 downto 0);
    signal count_inp1x_x1_834 : std_logic_vector(15 downto 0);
    signal count_inp1x_x1_900_delayed_1_0_915 : std_logic_vector(15 downto 0);
    signal count_inp1x_x1_at_entry_806 : std_logic_vector(15 downto 0);
    signal count_inp1x_x2_1317 : std_logic_vector(15 downto 0);
    signal count_inp2x_x0x_xph_1198 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_1049_delayed_3_0_1118 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_839 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_990_delayed_2_0_1032 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_at_entry_811 : std_logic_vector(15 downto 0);
    signal count_inp2x_x2_1343 : std_logic_vector(15 downto 0);
    signal exitcond1_1653 : std_logic_vector(0 downto 0);
    signal exitcond2_530 : std_logic_vector(0 downto 0);
    signal exitcond_752 : std_logic_vector(0 downto 0);
    signal forx_xbody169_forx_xend223x_xloopexit_taken_755 : std_logic_vector(0 downto 0);
    signal forx_xbody_forx_xcond163x_xpreheaderx_xloopexit_taken_533 : std_logic_vector(0 downto 0);
    signal iNsTr_19_346 : std_logic_vector(63 downto 0);
    signal iNsTr_33_568 : std_logic_vector(63 downto 0);
    signal iNsTr_81_1510 : std_logic_vector(63 downto 0);
    signal idxprom240_871 : std_logic_vector(63 downto 0);
    signal idxprom244_894 : std_logic_vector(63 downto 0);
    signal idxprom268_1074 : std_logic_vector(63 downto 0);
    signal idxprom272_1097 : std_logic_vector(63 downto 0);
    signal ifx_xend297_whilex_xend_taken_1355 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_950 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_968_delayed_1_0_1003 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_975_delayed_1_0_1012 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_980_delayed_1_0_1020 : std_logic_vector(0 downto 0);
    signal ifx_xend_ifx_xend297_taken_1026 : std_logic_vector(0 downto 0);
    signal ifx_xend_landx_xlhsx_xtrue_taken_1017 : std_logic_vector(0 downto 0);
    signal ifx_xthen266_exec_guard_1025_delayed_7_0_1084 : std_logic_vector(0 downto 0);
    signal ifx_xthen266_exec_guard_1042_delayed_13_0_1107 : std_logic_vector(0 downto 0);
    signal ifx_xthen266_exec_guard_1066 : std_logic_vector(0 downto 0);
    signal ifx_xthen266_landx_xlhsx_xtrue288_taken_1148 : std_logic_vector(0 downto 0);
    signal ifx_xthen296_exec_guard_1232 : std_logic_vector(0 downto 0);
    signal ifx_xthen296_ifx_xend297_taken_1235 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_863 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_876_delayed_7_0_881 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_893_delayed_13_0_904 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend_taken_945 : std_logic_vector(0 downto 0);
    signal inc247_922 : std_logic_vector(15 downto 0);
    signal inc249_932 : std_logic_vector(15 downto 0);
    signal inc251_942 : std_logic_vector(15 downto 0);
    signal inc275_1125 : std_logic_vector(15 downto 0);
    signal inc277_1135 : std_logic_vector(15 downto 0);
    signal inc279_1145 : std_logic_vector(15 downto 0);
    signal indvar476_592 : std_logic_vector(63 downto 0);
    signal indvar476_at_entry_584 : std_logic_vector(63 downto 0);
    signal indvar488_370 : std_logic_vector(63 downto 0);
    signal indvar488_at_entry_362 : std_logic_vector(63 downto 0);
    signal indvar_1526 : std_logic_vector(63 downto 0);
    signal indvarx_xnext477_747 : std_logic_vector(63 downto 0);
    signal indvarx_xnext489_525 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1648 : std_logic_vector(63 downto 0);
    signal landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1206 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1215 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1223 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue288_exec_guard_1153 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue288_ifx_xend297_taken_1229 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue288_ifx_xthen296_taken_1220 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_1029 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1040 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_ifx_xthen266_taken_1054 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_landx_xlhsx_xtrue288_taken_1063 : std_logic_vector(0 downto 0);
    signal mul105_280 : std_logic_vector(31 downto 0);
    signal mul111_291 : std_logic_vector(31 downto 0);
    signal mul85_259 : std_logic_vector(31 downto 0);
    signal mul91_264 : std_logic_vector(31 downto 0);
    signal mul98_269 : std_logic_vector(31 downto 0);
    signal mul_254 : std_logic_vector(31 downto 0);
    signal ptr_deref_1088_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1088_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1113_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1113_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1543_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_517_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_517_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_517_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_517_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_517_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_517_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_739_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_739_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_739_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_739_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_739_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_739_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_885_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_885_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_885_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_885_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_885_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_910_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_910_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_910_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_910_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_910_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_910_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl119_395 : std_logic_vector(63 downto 0);
    signal shl125_413 : std_logic_vector(63 downto 0);
    signal shl131_431 : std_logic_vector(63 downto 0);
    signal shl137_449 : std_logic_vector(63 downto 0);
    signal shl143_467 : std_logic_vector(63 downto 0);
    signal shl149_485 : std_logic_vector(63 downto 0);
    signal shl155_503 : std_logic_vector(63 downto 0);
    signal shl175_617 : std_logic_vector(63 downto 0);
    signal shl181_635 : std_logic_vector(63 downto 0);
    signal shl187_653 : std_logic_vector(63 downto 0);
    signal shl18_87 : std_logic_vector(31 downto 0);
    signal shl193_671 : std_logic_vector(63 downto 0);
    signal shl199_689 : std_logic_vector(63 downto 0);
    signal shl205_707 : std_logic_vector(63 downto 0);
    signal shl211_725 : std_logic_vector(63 downto 0);
    signal shl27_112 : std_logic_vector(31 downto 0);
    signal shl36_137 : std_logic_vector(31 downto 0);
    signal shl45_162 : std_logic_vector(31 downto 0);
    signal shl54_187 : std_logic_vector(31 downto 0);
    signal shl63_212 : std_logic_vector(31 downto 0);
    signal shl72_237 : std_logic_vector(31 downto 0);
    signal shl9_62 : std_logic_vector(31 downto 0);
    signal shl_37 : std_logic_vector(31 downto 0);
    signal shr236454_775 : std_logic_vector(31 downto 0);
    signal shr263458_781 : std_logic_vector(31 downto 0);
    signal shr301_787 : std_logic_vector(31 downto 0);
    signal shr317_1392 : std_logic_vector(63 downto 0);
    signal shr323_1402 : std_logic_vector(63 downto 0);
    signal shr329_1412 : std_logic_vector(63 downto 0);
    signal shr335_1422 : std_logic_vector(63 downto 0);
    signal shr341_1432 : std_logic_vector(63 downto 0);
    signal shr347_1442 : std_logic_vector(63 downto 0);
    signal shr353_1452 : std_logic_vector(63 downto 0);
    signal shr393_1554 : std_logic_vector(63 downto 0);
    signal shr399_1564 : std_logic_vector(63 downto 0);
    signal shr405_1574 : std_logic_vector(63 downto 0);
    signal shr411_1584 : std_logic_vector(63 downto 0);
    signal shr417_1594 : std_logic_vector(63 downto 0);
    signal shr423_1604 : std_logic_vector(63 downto 0);
    signal shr429_1614 : std_logic_vector(63 downto 0);
    signal sub_1382 : std_logic_vector(63 downto 0);
    signal tmp242_886 : std_logic_vector(63 downto 0);
    signal tmp270_1089 : std_logic_vector(63 downto 0);
    signal tmp386_1544 : std_logic_vector(63 downto 0);
    signal tmp471x_xop_1506 : std_logic_vector(31 downto 0);
    signal tmp472_1500 : std_logic_vector(0 downto 0);
    signal tmp475_1523 : std_logic_vector(63 downto 0);
    signal tmp480_546 : std_logic_vector(31 downto 0);
    signal tmp481_552 : std_logic_vector(31 downto 0);
    signal tmp481x_xop_564 : std_logic_vector(31 downto 0);
    signal tmp482_558 : std_logic_vector(0 downto 0);
    signal tmp486_581 : std_logic_vector(63 downto 0);
    signal tmp492_324 : std_logic_vector(31 downto 0);
    signal tmp493_330 : std_logic_vector(31 downto 0);
    signal tmp493x_xop_342 : std_logic_vector(31 downto 0);
    signal tmp494_336 : std_logic_vector(0 downto 0);
    signal tmp498_359 : std_logic_vector(63 downto 0);
    signal type_cast_1082_1082_delayed_2_0_1157 : std_logic_vector(15 downto 0);
    signal type_cast_1094_1094_delayed_3_0_1172 : std_logic_vector(15 downto 0);
    signal type_cast_1106_1106_delayed_3_0_1187 : std_logic_vector(15 downto 0);
    signal type_cast_110_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1123_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1143_1143_delayed_1_0_1239 : std_logic_vector(15 downto 0);
    signal type_cast_1143_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1146_1146_delayed_1_0_1243 : std_logic_vector(15 downto 0);
    signal type_cast_1149_1149_delayed_2_0_1247 : std_logic_vector(15 downto 0);
    signal type_cast_1159_1159_delayed_1_0_1267 : std_logic_vector(15 downto 0);
    signal type_cast_1161_wire : std_logic_vector(15 downto 0);
    signal type_cast_1162_1162_delayed_1_0_1271 : std_logic_vector(15 downto 0);
    signal type_cast_1165_1165_delayed_1_0_1275 : std_logic_vector(15 downto 0);
    signal type_cast_1165_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1176_wire : std_logic_vector(15 downto 0);
    signal type_cast_1179_1179_delayed_3_0_1295 : std_logic_vector(15 downto 0);
    signal type_cast_1180_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1182_1182_delayed_1_0_1299 : std_logic_vector(15 downto 0);
    signal type_cast_1191_wire : std_logic_vector(15 downto 0);
    signal type_cast_1195_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1196_1196_delayed_1_0_1321 : std_logic_vector(15 downto 0);
    signal type_cast_1199_1199_delayed_2_0_1325 : std_logic_vector(15 downto 0);
    signal type_cast_1252_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1280_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1304_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1311_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1330_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1337_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_135_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1367_wire : std_logic_vector(63 downto 0);
    signal type_cast_1375_wire : std_logic_vector(63 downto 0);
    signal type_cast_1390_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1400_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1410_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1440_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1450_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1485_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1498_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1504_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1514_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1521_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1530_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1532_wire : std_logic_vector(63 downto 0);
    signal type_cast_1552_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1562_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1572_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1582_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1592_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1602_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_160_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1612_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1646_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_210_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_235_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_273_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_284_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_295_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_310_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_328_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_334_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_340_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_357_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_35_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_373_wire : std_logic_vector(63 downto 0);
    signal type_cast_393_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_411_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_429_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_465_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_483_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_501_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_523_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_550_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_556_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_562_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_572_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_579_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_595_wire : std_logic_vector(63 downto 0);
    signal type_cast_60_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_615_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_633_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_651_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_669_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_687_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_705_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_723_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_745_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_779_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_785_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_822_wire : std_logic_vector(15 downto 0);
    signal type_cast_827_wire : std_logic_vector(15 downto 0);
    signal type_cast_832_wire : std_logic_vector(15 downto 0);
    signal type_cast_837_wire : std_logic_vector(15 downto 0);
    signal type_cast_842_wire : std_logic_vector(15 downto 0);
    signal type_cast_85_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_930_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_933_933_delayed_1_0_954 : std_logic_vector(15 downto 0);
    signal type_cast_940_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_945_945_delayed_1_0_969 : std_logic_vector(15 downto 0);
    signal type_cast_957_957_delayed_1_0_984 : std_logic_vector(15 downto 0);
    signal type_cast_958_wire : std_logic_vector(15 downto 0);
    signal type_cast_962_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_973_wire : std_logic_vector(15 downto 0);
    signal type_cast_977_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_988_wire : std_logic_vector(15 downto 0);
    signal type_cast_992_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_ifx_xend_taken_860 : std_logic_vector(0 downto 0);
    signal whilex_xbody_ifx_xthen_taken_856 : std_logic_vector(0 downto 0);
    signal xx_xop500_574 : std_logic_vector(63 downto 0);
    signal xx_xop501_352 : std_logic_vector(63 downto 0);
    signal xx_xop_1516 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    add_inp1x_x1_at_entry_796 <= "0000000000000000";
    add_inp2x_x1_at_entry_801 <= "0000000000000000";
    add_outx_x1_at_entry_790 <= "0000000000000000";
    array_obj_ref_1079_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1079_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1079_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1079_resized_base_address <= "00000000000000";
    array_obj_ref_1102_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1102_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1102_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1102_resized_base_address <= "00000000000000";
    array_obj_ref_1538_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1538_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1538_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1538_resized_base_address <= "00000000000000";
    array_obj_ref_380_constant_part_of_offset <= "00000000000000";
    array_obj_ref_380_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_380_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_380_resized_base_address <= "00000000000000";
    array_obj_ref_602_constant_part_of_offset <= "00000000000000";
    array_obj_ref_602_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_602_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_602_resized_base_address <= "00000000000000";
    array_obj_ref_876_constant_part_of_offset <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_876_resized_base_address <= "00000000000000";
    array_obj_ref_899_constant_part_of_offset <= "00000000000000";
    array_obj_ref_899_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_899_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_899_resized_base_address <= "00000000000000";
    count_inp1x_x1_at_entry_806 <= "0000000000000000";
    count_inp2x_x1_at_entry_811 <= "0000000000000000";
    indvar476_at_entry_584 <= "0000000000000000000000000000000000000000000000000000000000000000";
    indvar488_at_entry_362 <= "0000000000000000000000000000000000000000000000000000000000000000";
    ptr_deref_1088_word_offset_0 <= "00000000000000";
    ptr_deref_1113_word_offset_0 <= "00000000000000";
    ptr_deref_1543_word_offset_0 <= "00000000000000";
    ptr_deref_517_word_offset_0 <= "00000000000000";
    ptr_deref_739_word_offset_0 <= "00000000000000";
    ptr_deref_885_word_offset_0 <= "00000000000000";
    ptr_deref_910_word_offset_0 <= "00000000000000";
    type_cast_110_wire_constant <= "00000000000000000000000000001000";
    type_cast_1123_wire_constant <= "0000000000000001";
    type_cast_1133_wire_constant <= "0000000000000001";
    type_cast_1143_wire_constant <= "0000000000000001";
    type_cast_1165_wire_constant <= "0000000000000000";
    type_cast_1180_wire_constant <= "0000000000000000";
    type_cast_1195_wire_constant <= "0000000000000000";
    type_cast_1252_wire_constant <= "0000000000000000";
    type_cast_1280_wire_constant <= "0000000000000000";
    type_cast_1304_wire_constant <= "0000000000000000";
    type_cast_1311_wire_constant <= "0000000000000000";
    type_cast_1330_wire_constant <= "0000000000000000";
    type_cast_1337_wire_constant <= "0000000000000000";
    type_cast_135_wire_constant <= "00000000000000000000000000001000";
    type_cast_1390_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1400_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1410_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1420_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1430_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1440_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1450_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1485_wire_constant <= "00000000000000000000000000000111";
    type_cast_1498_wire_constant <= "00000000000000000000000000000001";
    type_cast_1504_wire_constant <= "11111111111111111111111111111111";
    type_cast_1514_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1521_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1530_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1552_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1562_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1572_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1582_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1592_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1602_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_160_wire_constant <= "00000000000000000000000000001000";
    type_cast_1612_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1646_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_185_wire_constant <= "00000000000000000000000000001000";
    type_cast_210_wire_constant <= "00000000000000000000000000001000";
    type_cast_235_wire_constant <= "00000000000000000000000000001000";
    type_cast_273_wire_constant <= "00000000000000001111111111111111";
    type_cast_284_wire_constant <= "00000000000000001111111111111111";
    type_cast_295_wire_constant <= "00000000000000000000000000000111";
    type_cast_310_wire_constant <= "00000000000000000000000000000111";
    type_cast_328_wire_constant <= "00000000000000000000000000000011";
    type_cast_334_wire_constant <= "00000000000000000000000000000001";
    type_cast_340_wire_constant <= "11111111111111111111111111111111";
    type_cast_350_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_357_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_35_wire_constant <= "00000000000000000000000000001000";
    type_cast_393_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_411_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_429_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_447_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_465_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_483_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_501_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_523_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_550_wire_constant <= "00000000000000000000000000000011";
    type_cast_556_wire_constant <= "00000000000000000000000000000001";
    type_cast_562_wire_constant <= "11111111111111111111111111111111";
    type_cast_572_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_579_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_60_wire_constant <= "00000000000000000000000000001000";
    type_cast_615_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_633_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_651_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_669_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_687_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_705_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_723_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_745_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_773_wire_constant <= "00000000000000000000000000000011";
    type_cast_779_wire_constant <= "00000000000000000000000000000011";
    type_cast_785_wire_constant <= "00000000000000000000000000000011";
    type_cast_85_wire_constant <= "00000000000000000000000000001000";
    type_cast_920_wire_constant <= "0000000000000001";
    type_cast_930_wire_constant <= "0000000000000001";
    type_cast_940_wire_constant <= "0000000000000001";
    type_cast_962_wire_constant <= "0000000000000000";
    type_cast_977_wire_constant <= "0000000000000000";
    type_cast_992_wire_constant <= "0000000000000000";
    phi_stmt_1526: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1530_wire_constant & type_cast_1532_wire;
      req <= phi_stmt_1526_req_0 & phi_stmt_1526_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1526",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1526_ack_0,
          idata => idata,
          odata => indvar_1526,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1526
    phi_stmt_370: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_373_wire & indvar488_at_entry_362;
      req <= phi_stmt_370_req_0 & phi_stmt_370_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_370",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_370_ack_0,
          idata => idata,
          odata => indvar488_370,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_370
    phi_stmt_592: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_595_wire & indvar476_at_entry_584;
      req <= phi_stmt_592_req_0 & phi_stmt_592_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_592",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_592_ack_0,
          idata => idata,
          odata => indvar476_592,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_592
    phi_stmt_819: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_822_wire & add_outx_x1_at_entry_790;
      req <= phi_stmt_819_req_0 & phi_stmt_819_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_819",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_819_ack_0,
          idata => idata,
          odata => add_outx_x1_819,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_819
    phi_stmt_824: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_827_wire & add_inp1x_x1_at_entry_796;
      req <= phi_stmt_824_req_0 & phi_stmt_824_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_824",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_824_ack_0,
          idata => idata,
          odata => add_inp1x_x1_824,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_824
    phi_stmt_829: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_832_wire & add_inp2x_x1_at_entry_801;
      req <= phi_stmt_829_req_0 & phi_stmt_829_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_829",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_829_ack_0,
          idata => idata,
          odata => add_inp2x_x1_829,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_829
    phi_stmt_834: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_837_wire & count_inp1x_x1_at_entry_806;
      req <= phi_stmt_834_req_0 & phi_stmt_834_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_834",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_834_ack_0,
          idata => idata,
          odata => count_inp1x_x1_834,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_834
    phi_stmt_839: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_842_wire & count_inp2x_x1_at_entry_811;
      req <= phi_stmt_839_req_0 & phi_stmt_839_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_839",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_839_ack_0,
          idata => idata,
          odata => count_inp2x_x1_839,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_839
    -- flow-through select operator MUX_1166_inst
    MUX_1166_wire <= type_cast_1082_1082_delayed_2_0_1157 when (landx_xlhsx_xtrue_landx_xlhsx_xtrue288_taken_1063(0) /=  '0') else type_cast_1165_wire_constant;
    -- flow-through select operator MUX_1167_inst
    add_outx_x2x_xph_1168 <= type_cast_1161_wire when (ifx_xthen266_landx_xlhsx_xtrue288_taken_1148(0) /=  '0') else MUX_1166_wire;
    -- flow-through select operator MUX_1181_inst
    MUX_1181_wire <= type_cast_1094_1094_delayed_3_0_1172 when (landx_xlhsx_xtrue_landx_xlhsx_xtrue288_taken_1063(0) /=  '0') else type_cast_1180_wire_constant;
    -- flow-through select operator MUX_1182_inst
    add_inp2x_x0x_xph_1183 <= type_cast_1176_wire when (ifx_xthen266_landx_xlhsx_xtrue288_taken_1148(0) /=  '0') else MUX_1181_wire;
    -- flow-through select operator MUX_1196_inst
    MUX_1196_wire <= type_cast_1106_1106_delayed_3_0_1187 when (landx_xlhsx_xtrue_landx_xlhsx_xtrue288_taken_1063(0) /=  '0') else type_cast_1195_wire_constant;
    -- flow-through select operator MUX_1197_inst
    count_inp2x_x0x_xph_1198 <= type_cast_1191_wire when (ifx_xthen266_landx_xlhsx_xtrue288_taken_1148(0) /=  '0') else MUX_1196_wire;
    MUX_1253_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1253_inst_req_0;
      MUX_1253_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1253_inst_req_1;
      MUX_1253_inst_ack_1<= update_ack(0);
      MUX_1253_inst: SelectSplitProtocol generic map(name => "MUX_1253_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1149_1149_delayed_2_0_1247, y => type_cast_1252_wire_constant, sel => ifx_xend_ifx_xend297_taken_1026, z => MUX_1152_1152_delayed_2_0_1254, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1261_inst
    MUX_1261_wire <= type_cast_1146_1146_delayed_1_0_1243 when (landx_xlhsx_xtrue288_ifx_xend297_taken_1229(0) /=  '0') else MUX_1152_1152_delayed_2_0_1254;
    -- flow-through select operator MUX_1262_inst
    add_inp2x_x0504_1263 <= type_cast_1143_1143_delayed_1_0_1239 when (ifx_xthen296_ifx_xend297_taken_1235(0) /=  '0') else MUX_1261_wire;
    MUX_1281_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1281_inst_req_0;
      MUX_1281_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1281_inst_req_1;
      MUX_1281_inst_ack_1<= update_ack(0);
      MUX_1281_inst: SelectSplitProtocol generic map(name => "MUX_1281_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1165_1165_delayed_1_0_1275, y => type_cast_1280_wire_constant, sel => ifx_xend_ifx_xend297_taken_1026, z => MUX_1168_1168_delayed_2_0_1282, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1289_inst
    MUX_1289_wire <= type_cast_1162_1162_delayed_1_0_1271 when (landx_xlhsx_xtrue288_ifx_xend297_taken_1229(0) /=  '0') else MUX_1168_1168_delayed_2_0_1282;
    -- flow-through select operator MUX_1290_inst
    add_outx_x2502_1291 <= type_cast_1159_1159_delayed_1_0_1267 when (ifx_xthen296_ifx_xend297_taken_1235(0) /=  '0') else MUX_1289_wire;
    MUX_1305_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1305_inst_req_0;
      MUX_1305_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1305_inst_req_1;
      MUX_1305_inst_ack_1<= update_ack(0);
      MUX_1305_inst: SelectSplitProtocol generic map(name => "MUX_1305_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1182_1182_delayed_1_0_1299, y => type_cast_1304_wire_constant, sel => ifx_xend_ifx_xend297_taken_1026, z => MUX_1185_1185_delayed_2_0_1306, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1315_inst
    MUX_1315_wire <= type_cast_1179_1179_delayed_3_0_1295 when (landx_xlhsx_xtrue288_ifx_xend297_taken_1229(0) /=  '0') else MUX_1185_1185_delayed_2_0_1306;
    -- flow-through select operator MUX_1316_inst
    count_inp1x_x2_1317 <= type_cast_1311_wire_constant when (ifx_xthen296_ifx_xend297_taken_1235(0) /=  '0') else MUX_1315_wire;
    MUX_1331_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1331_inst_req_0;
      MUX_1331_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1331_inst_req_1;
      MUX_1331_inst_ack_1<= update_ack(0);
      MUX_1331_inst: SelectSplitProtocol generic map(name => "MUX_1331_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1199_1199_delayed_2_0_1325, y => type_cast_1330_wire_constant, sel => ifx_xend_ifx_xend297_taken_1026, z => MUX_1202_1202_delayed_2_0_1332, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1341_inst
    MUX_1341_wire <= type_cast_1196_1196_delayed_1_0_1321 when (landx_xlhsx_xtrue288_ifx_xend297_taken_1229(0) /=  '0') else MUX_1202_1202_delayed_2_0_1332;
    -- flow-through select operator MUX_1342_inst
    count_inp2x_x2_1343 <= type_cast_1337_wire_constant when (ifx_xthen296_ifx_xend297_taken_1235(0) /=  '0') else MUX_1341_wire;
    -- flow-through select operator MUX_1522_inst
    tmp475_1523 <= xx_xop_1516 when (tmp472_1500(0) /=  '0') else type_cast_1521_wire_constant;
    -- flow-through select operator MUX_358_inst
    tmp498_359 <= xx_xop501_352 when (tmp494_336(0) /=  '0') else type_cast_357_wire_constant;
    -- flow-through select operator MUX_580_inst
    tmp486_581 <= xx_xop500_574 when (tmp482_558(0) /=  '0') else type_cast_579_wire_constant;
    -- flow-through select operator MUX_963_inst
    MUX_963_wire <= type_cast_933_933_delayed_1_0_954 when (whilex_xbody_ifx_xend_taken_860(0) /=  '0') else type_cast_962_wire_constant;
    -- flow-through select operator MUX_964_inst
    add_outx_x0_965 <= type_cast_958_wire when (ifx_xthen_ifx_xend_taken_945(0) /=  '0') else MUX_963_wire;
    -- flow-through select operator MUX_978_inst
    MUX_978_wire <= type_cast_945_945_delayed_1_0_969 when (whilex_xbody_ifx_xend_taken_860(0) /=  '0') else type_cast_977_wire_constant;
    -- flow-through select operator MUX_979_inst
    add_inp1x_x0_980 <= type_cast_973_wire when (ifx_xthen_ifx_xend_taken_945(0) /=  '0') else MUX_978_wire;
    -- flow-through select operator MUX_993_inst
    MUX_993_wire <= type_cast_957_957_delayed_1_0_984 when (whilex_xbody_ifx_xend_taken_860(0) /=  '0') else type_cast_992_wire_constant;
    -- flow-through select operator MUX_994_inst
    count_inp1x_x0_995 <= type_cast_988_wire when (ifx_xthen_ifx_xend_taken_945(0) /=  '0') else MUX_993_wire;
    W_add_inp1x_x1_866_delayed_1_0_864_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp1x_x1_866_delayed_1_0_864_inst_req_0;
      W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp1x_x1_866_delayed_1_0_864_inst_req_1;
      W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_1<= rack(0);
      W_add_inp1x_x1_866_delayed_1_0_864_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp1x_x1_866_delayed_1_0_864_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp1x_x1_866_delayed_1_0_866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_inp1x_x1_907_delayed_1_0_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp1x_x1_907_delayed_1_0_923_inst_req_0;
      W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp1x_x1_907_delayed_1_0_923_inst_req_1;
      W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_1<= rack(0);
      W_add_inp1x_x1_907_delayed_1_0_923_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp1x_x1_907_delayed_1_0_923_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp1x_x1_907_delayed_1_0_925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_inp2x_x1_1015_delayed_3_0_1067_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_0;
      W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_1;
      W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_1<= rack(0);
      W_add_inp2x_x1_1015_delayed_3_0_1067_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp2x_x1_1015_delayed_3_0_1067_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp2x_x1_1015_delayed_3_0_1069,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_inp2x_x1_1056_delayed_3_0_1126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_0;
      W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_1;
      W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_1<= rack(0);
      W_add_inp2x_x1_1056_delayed_3_0_1126_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp2x_x1_1056_delayed_3_0_1126_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp2x_x1_1056_delayed_3_0_1128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x0_1032_delayed_2_0_1090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x0_1032_delayed_2_0_1090_inst_req_0;
      W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x0_1032_delayed_2_0_1090_inst_req_1;
      W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_1<= rack(0);
      W_add_outx_x0_1032_delayed_2_0_1090_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x0_1032_delayed_2_0_1090_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x0_1032_delayed_2_0_1092,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x0_1063_delayed_2_0_1136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x0_1063_delayed_2_0_1136_inst_req_0;
      W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x0_1063_delayed_2_0_1136_inst_req_1;
      W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_1<= rack(0);
      W_add_outx_x0_1063_delayed_2_0_1136_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x0_1063_delayed_2_0_1136_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x0_1063_delayed_2_0_1138,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x1_883_delayed_1_0_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x1_883_delayed_1_0_887_inst_req_0;
      W_add_outx_x1_883_delayed_1_0_887_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x1_883_delayed_1_0_887_inst_req_1;
      W_add_outx_x1_883_delayed_1_0_887_inst_ack_1<= rack(0);
      W_add_outx_x1_883_delayed_1_0_887_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x1_883_delayed_1_0_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x1_883_delayed_1_0_889,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x1_914_delayed_1_0_933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x1_914_delayed_1_0_933_inst_req_0;
      W_add_outx_x1_914_delayed_1_0_933_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x1_914_delayed_1_0_933_inst_req_1;
      W_add_outx_x1_914_delayed_1_0_933_inst_ack_1<= rack(0);
      W_add_outx_x1_914_delayed_1_0_933_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x1_914_delayed_1_0_933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x1_914_delayed_1_0_935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx245_894_delayed_6_0_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx245_894_delayed_6_0_905_inst_req_0;
      W_arrayidx245_894_delayed_6_0_905_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx245_894_delayed_6_0_905_inst_req_1;
      W_arrayidx245_894_delayed_6_0_905_inst_ack_1<= rack(0);
      W_arrayidx245_894_delayed_6_0_905_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx245_894_delayed_6_0_905_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx245_901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx245_894_delayed_6_0_907,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx273_1043_delayed_6_0_1108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx273_1043_delayed_6_0_1108_inst_req_0;
      W_arrayidx273_1043_delayed_6_0_1108_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx273_1043_delayed_6_0_1108_inst_req_1;
      W_arrayidx273_1043_delayed_6_0_1108_inst_ack_1<= rack(0);
      W_arrayidx273_1043_delayed_6_0_1108_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx273_1043_delayed_6_0_1108_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx273_1104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx273_1043_delayed_6_0_1110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_inp1x_x1_900_delayed_1_0_913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_inp1x_x1_900_delayed_1_0_913_inst_req_0;
      W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_0<= wack(0);
      rreq(0) <= W_count_inp1x_x1_900_delayed_1_0_913_inst_req_1;
      W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_1<= rack(0);
      W_count_inp1x_x1_900_delayed_1_0_913_inst : InterlockBuffer generic map ( -- 
        name => "W_count_inp1x_x1_900_delayed_1_0_913_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x1_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_inp1x_x1_900_delayed_1_0_915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_inp2x_x1_1049_delayed_3_0_1116_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_0;
      W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_0<= wack(0);
      rreq(0) <= W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_1;
      W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_1<= rack(0);
      W_count_inp2x_x1_1049_delayed_3_0_1116_inst : InterlockBuffer generic map ( -- 
        name => "W_count_inp2x_x1_1049_delayed_3_0_1116_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_inp2x_x1_1049_delayed_3_0_1118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_inp2x_x1_990_delayed_2_0_1030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_0;
      W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_0<= wack(0);
      rreq(0) <= W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_1;
      W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_1<= rack(0);
      W_count_inp2x_x1_990_delayed_2_0_1030_inst : InterlockBuffer generic map ( -- 
        name => "W_count_inp2x_x1_990_delayed_2_0_1030_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_inp2x_x1_990_delayed_2_0_1032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_forx_xbody169_forx_xend223x_xloopexit_taken_753_inst
    process(exitcond_752) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := exitcond_752(0 downto 0);
      forx_xbody169_forx_xend223x_xloopexit_taken_755 <= tmp_var; -- 
    end process;
    -- interlock W_forx_xbody_forx_xcond163x_xpreheaderx_xloopexit_taken_531_inst
    process(exitcond2_530) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := exitcond2_530(0 downto 0);
      forx_xbody_forx_xcond163x_xpreheaderx_xloopexit_taken_533 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xend297_whilex_xend_taken_1353_inst
    process(cmp302_1352) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp302_1352(0 downto 0);
      ifx_xend297_whilex_xend_taken_1355 <= tmp_var; -- 
    end process;
    W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_0;
      W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_1;
      W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_968_delayed_1_0_1003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_0;
      W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_1;
      W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_975_delayed_1_0_1012,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_0;
      W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_1;
      W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_980_delayed_1_0_1020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_req_0;
      W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_req_1;
      W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst_ack_1<= rack(0);
      W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen266_exec_guard_1025_delayed_7_0_1082_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen266_exec_guard_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen266_exec_guard_1025_delayed_7_0_1084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_req_0;
      W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_req_1;
      W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst_ack_1<= rack(0);
      W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen266_exec_guard_1042_delayed_13_0_1105_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen266_exec_guard_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen266_exec_guard_1042_delayed_13_0_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen266_exec_guard_1064_inst
    process(landx_xlhsx_xtrue_ifx_xthen266_taken_1054) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := landx_xlhsx_xtrue_ifx_xthen266_taken_1054(0 downto 0);
      ifx_xthen266_exec_guard_1066 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen266_landx_xlhsx_xtrue288_taken_1146_inst
    process(ifx_xthen266_exec_guard_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen266_exec_guard_1066(0 downto 0);
      ifx_xthen266_landx_xlhsx_xtrue288_taken_1148 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen296_exec_guard_1230_inst
    process(landx_xlhsx_xtrue288_ifx_xthen296_taken_1220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := landx_xlhsx_xtrue288_ifx_xthen296_taken_1220(0 downto 0);
      ifx_xthen296_exec_guard_1232 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen296_ifx_xend297_taken_1233_inst
    process(ifx_xthen296_exec_guard_1232) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen296_exec_guard_1232(0 downto 0);
      ifx_xthen296_ifx_xend297_taken_1235 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen_exec_guard_861_inst
    process(whilex_xbody_ifx_xthen_taken_856) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xthen_taken_856(0 downto 0);
      ifx_xthen_exec_guard_863 <= tmp_var; -- 
    end process;
    W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_0;
      W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_1;
      W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_1<= rack(0);
      W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_exec_guard_863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_exec_guard_876_delayed_7_0_881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_0;
      W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_1;
      W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_1<= rack(0);
      W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_exec_guard_863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_exec_guard_893_delayed_13_0_904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen_ifx_xend_taken_943_inst
    process(ifx_xthen_exec_guard_863) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen_exec_guard_863(0 downto 0);
      ifx_xthen_ifx_xend_taken_945 <= tmp_var; -- 
    end process;
    W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_req_0;
      W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_req_1;
      W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1204_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue288_exec_guard_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue288_exec_guard_1117_delayed_1_0_1206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_req_0;
      W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_req_1;
      W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1213_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue288_exec_guard_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_req_0;
      W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_req_1;
      W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1221_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue288_exec_guard_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_0;
      W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_1;
      W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue_exec_guard_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_0;
      W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_1;
      W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue_exec_guard_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_landx_xlhsx_xtrue_exec_guard_1027_inst
    process(ifx_xend_landx_xlhsx_xtrue_taken_1017) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xend_landx_xlhsx_xtrue_taken_1017(0 downto 0);
      landx_xlhsx_xtrue_exec_guard_1029 <= tmp_var; -- 
    end process;
    W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_0;
      W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_1;
      W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue_exec_guard_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1040,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_ifx_xthen_taken_854_inst
    process(cmp237_853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp237_853(0 downto 0);
      whilex_xbody_ifx_xthen_taken_856 <= tmp_var; -- 
    end process;
    addr_of_1080_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1080_final_reg_req_0;
      addr_of_1080_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1080_final_reg_req_1;
      addr_of_1080_final_reg_ack_1<= rack(0);
      addr_of_1080_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1080_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1079_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_1081,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1103_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1103_final_reg_req_0;
      addr_of_1103_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1103_final_reg_req_1;
      addr_of_1103_final_reg_ack_1<= rack(0);
      addr_of_1103_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1103_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1102_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx273_1104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1539_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1539_final_reg_req_0;
      addr_of_1539_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1539_final_reg_req_1;
      addr_of_1539_final_reg_ack_1<= rack(0);
      addr_of_1539_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1539_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1538_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx385_1540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_381_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_381_final_reg_req_0;
      addr_of_381_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_381_final_reg_req_1;
      addr_of_381_final_reg_ack_1<= rack(0);
      addr_of_381_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_381_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_380_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_603_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_603_final_reg_req_0;
      addr_of_603_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_603_final_reg_req_1;
      addr_of_603_final_reg_ack_1<= rack(0);
      addr_of_603_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_603_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_602_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx219_604,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_877_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_877_final_reg_req_0;
      addr_of_877_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_877_final_reg_req_1;
      addr_of_877_final_reg_ack_1<= rack(0);
      addr_of_877_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_877_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_876_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx241_878,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_900_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_900_final_reg_req_0;
      addr_of_900_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_900_final_reg_req_1;
      addr_of_900_final_reg_ack_1<= rack(0);
      addr_of_900_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_900_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_899_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx245_901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1036_inst_req_0;
      type_cast_1036_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1036_inst_req_1;
      type_cast_1036_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  landx_xlhsx_xtrue_exec_guard_1029(0);
      type_cast_1036_inst_gI: SplitGuardInterface generic map(name => "type_cast_1036_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1036_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1036_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_990_delayed_2_0_1032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv260_1037,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_105_inst_req_0;
      type_cast_105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_105_inst_req_1;
      type_cast_105_inst_ack_1<= rack(0);
      type_cast_105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1073_inst_req_0;
      type_cast_1073_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1073_inst_req_1;
      type_cast_1073_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen266_exec_guard_1066(0);
      type_cast_1073_inst_gI: SplitGuardInterface generic map(name => "type_cast_1073_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1073_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1073_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_1015_delayed_3_0_1069,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom268_1074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1096_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1096_inst_req_0;
      type_cast_1096_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1096_inst_req_1;
      type_cast_1096_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen266_exec_guard_1066(0);
      type_cast_1096_inst_gI: SplitGuardInterface generic map(name => "type_cast_1096_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1096_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1096_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_1032_delayed_2_0_1092,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom272_1097,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1156_inst_req_0;
      type_cast_1156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1156_inst_req_1;
      type_cast_1156_inst_ack_1<= rack(0);
      type_cast_1156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1156_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1082_1082_delayed_2_0_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1161_inst
    process(inc279_1145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc279_1145(15 downto 0);
      type_cast_1161_wire <= tmp_var; -- 
    end process;
    type_cast_1171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1171_inst_req_0;
      type_cast_1171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1171_inst_req_1;
      type_cast_1171_inst_ack_1<= rack(0);
      type_cast_1171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1171_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1094_1094_delayed_3_0_1172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1176_inst
    process(inc277_1135) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc277_1135(15 downto 0);
      type_cast_1176_wire <= tmp_var; -- 
    end process;
    type_cast_1186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1186_inst_req_0;
      type_cast_1186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1186_inst_req_1;
      type_cast_1186_inst_ack_1<= rack(0);
      type_cast_1186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1186_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1106_1106_delayed_3_0_1187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_118_inst_req_0;
      type_cast_118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_118_inst_req_1;
      type_cast_118_inst_ack_1<= rack(0);
      type_cast_118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1191_inst
    process(inc275_1125) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc275_1125(15 downto 0);
      type_cast_1191_wire <= tmp_var; -- 
    end process;
    type_cast_1202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1202_inst_req_0;
      type_cast_1202_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1202_inst_req_1;
      type_cast_1202_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  landx_xlhsx_xtrue288_exec_guard_1153(0);
      type_cast_1202_inst_gI: SplitGuardInterface generic map(name => "type_cast_1202_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1202_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x0x_xph_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv290_1203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x0x_xph_1183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1143_1143_delayed_1_0_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1242_inst_req_0;
      type_cast_1242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1242_inst_req_1;
      type_cast_1242_inst_ack_1<= rack(0);
      type_cast_1242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1242_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x0x_xph_1183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1146_1146_delayed_1_0_1243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1246_inst_req_0;
      type_cast_1246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1246_inst_req_1;
      type_cast_1246_inst_ack_1<= rack(0);
      type_cast_1246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1246_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1149_1149_delayed_2_0_1247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1266_inst_req_0;
      type_cast_1266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1266_inst_req_1;
      type_cast_1266_inst_ack_1<= rack(0);
      type_cast_1266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1266_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2x_xph_1168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1159_1159_delayed_1_0_1267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1270_inst_req_0;
      type_cast_1270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1270_inst_req_1;
      type_cast_1270_inst_ack_1<= rack(0);
      type_cast_1270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1270_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2x_xph_1168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1162_1162_delayed_1_0_1271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1274_inst_req_0;
      type_cast_1274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1274_inst_req_1;
      type_cast_1274_inst_ack_1<= rack(0);
      type_cast_1274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1165_1165_delayed_1_0_1275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1294_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1294_inst_req_0;
      type_cast_1294_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1294_inst_req_1;
      type_cast_1294_inst_ack_1<= rack(0);
      type_cast_1294_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1294_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x0_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1179_1179_delayed_3_0_1295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1298_inst_req_0;
      type_cast_1298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1298_inst_req_1;
      type_cast_1298_inst_ack_1<= rack(0);
      type_cast_1298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x0_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1182_1182_delayed_1_0_1299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_130_inst_req_0;
      type_cast_130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_130_inst_req_1;
      type_cast_130_inst_ack_1<= rack(0);
      type_cast_130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1320_inst_req_0;
      type_cast_1320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1320_inst_req_1;
      type_cast_1320_inst_ack_1<= rack(0);
      type_cast_1320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1320_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x0x_xph_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1196_1196_delayed_1_0_1321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1324_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1324_inst_req_0;
      type_cast_1324_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1324_inst_req_1;
      type_cast_1324_inst_ack_1<= rack(0);
      type_cast_1324_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1324_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1199_1199_delayed_2_0_1325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1346_inst_req_0;
      type_cast_1346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1346_inst_req_1;
      type_cast_1346_inst_ack_1<= rack(0);
      type_cast_1346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2502_1291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv299_1347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1368_inst_req_0;
      type_cast_1368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1368_inst_req_1;
      type_cast_1368_inst_ack_1<= rack(0);
      type_cast_1368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1367_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv226_1369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1376_inst_req_0;
      type_cast_1376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1376_inst_req_1;
      type_cast_1376_inst_ack_1<= rack(0);
      type_cast_1376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1375_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv308_1377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1385_inst_req_0;
      type_cast_1385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1385_inst_req_1;
      type_cast_1385_inst_ack_1<= rack(0);
      type_cast_1385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv314_1386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1395_inst_req_0;
      type_cast_1395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1395_inst_req_1;
      type_cast_1395_inst_ack_1<= rack(0);
      type_cast_1395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr317_1392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv320_1396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1405_inst_req_0;
      type_cast_1405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1405_inst_req_1;
      type_cast_1405_inst_ack_1<= rack(0);
      type_cast_1405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr323_1402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv326_1406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1415_inst_req_0;
      type_cast_1415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1415_inst_req_1;
      type_cast_1415_inst_ack_1<= rack(0);
      type_cast_1415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1415_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr329_1412,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv332_1416,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1425_inst_req_0;
      type_cast_1425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1425_inst_req_1;
      type_cast_1425_inst_ack_1<= rack(0);
      type_cast_1425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr335_1422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv338_1426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1435_inst_req_0;
      type_cast_1435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1435_inst_req_1;
      type_cast_1435_inst_ack_1<= rack(0);
      type_cast_1435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr341_1432,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv344_1436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_143_inst_req_0;
      type_cast_143_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_143_inst_req_1;
      type_cast_143_inst_ack_1<= rack(0);
      type_cast_143_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_140,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_144,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1445_inst_req_0;
      type_cast_1445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1445_inst_req_1;
      type_cast_1445_inst_ack_1<= rack(0);
      type_cast_1445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr347_1442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv350_1446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1455_inst_req_0;
      type_cast_1455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1455_inst_req_1;
      type_cast_1455_inst_ack_1<= rack(0);
      type_cast_1455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr353_1452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv356_1456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1509_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1509_inst_req_0;
      type_cast_1509_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1509_inst_req_1;
      type_cast_1509_inst_ack_1<= rack(0);
      type_cast_1509_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1509_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp471x_xop_1506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_81_1510,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1532_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1532_inst_req_0;
      type_cast_1532_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1532_inst_req_1;
      type_cast_1532_inst_ack_1<= rack(0);
      type_cast_1532_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1532_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1532_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1547_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1547_inst_req_0;
      type_cast_1547_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1547_inst_req_1;
      type_cast_1547_inst_ack_1<= rack(0);
      type_cast_1547_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1547_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp386_1544,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv390_1548,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1557_inst_req_0;
      type_cast_1557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1557_inst_req_1;
      type_cast_1557_inst_ack_1<= rack(0);
      type_cast_1557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr393_1554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv396_1558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1567_inst_req_0;
      type_cast_1567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1567_inst_req_1;
      type_cast_1567_inst_ack_1<= rack(0);
      type_cast_1567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr399_1564,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv402_1568,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1577_inst_req_0;
      type_cast_1577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1577_inst_req_1;
      type_cast_1577_inst_ack_1<= rack(0);
      type_cast_1577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr405_1574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv408_1578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1587_inst_req_0;
      type_cast_1587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1587_inst_req_1;
      type_cast_1587_inst_ack_1<= rack(0);
      type_cast_1587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr411_1584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv414_1588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1597_inst_req_0;
      type_cast_1597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1597_inst_req_1;
      type_cast_1597_inst_ack_1<= rack(0);
      type_cast_1597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr417_1594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv420_1598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1607_inst_req_0;
      type_cast_1607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1607_inst_req_1;
      type_cast_1607_inst_ack_1<= rack(0);
      type_cast_1607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr423_1604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv426_1608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1617_inst_req_0;
      type_cast_1617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1617_inst_req_1;
      type_cast_1617_inst_ack_1<= rack(0);
      type_cast_1617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1617_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr429_1614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv432_1618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_168_inst_req_0;
      type_cast_168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_168_inst_req_1;
      type_cast_168_inst_ack_1<= rack(0);
      type_cast_168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_180_inst_req_0;
      type_cast_180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_180_inst_req_1;
      type_cast_180_inst_ack_1<= rack(0);
      type_cast_180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_193_inst_req_0;
      type_cast_193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_193_inst_req_1;
      type_cast_193_inst_ack_1<= rack(0);
      type_cast_193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_205_inst_req_0;
      type_cast_205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_205_inst_req_1;
      type_cast_205_inst_ack_1<= rack(0);
      type_cast_205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call59_202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_218_inst_req_0;
      type_cast_218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_218_inst_req_1;
      type_cast_218_inst_ack_1<= rack(0);
      type_cast_218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call64_215,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_230_inst_req_0;
      type_cast_230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_230_inst_req_1;
      type_cast_230_inst_ack_1<= rack(0);
      type_cast_230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_227,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_243_inst_req_0;
      type_cast_243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_243_inst_req_1;
      type_cast_243_inst_ack_1<= rack(0);
      type_cast_243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call73_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_30_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_30_inst_req_0;
      type_cast_30_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_30_inst_req_1;
      type_cast_30_inst_ack_1<= rack(0);
      type_cast_30_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_30_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_26,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_31,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp493x_xop_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_19_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_373_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_373_inst_req_0;
      type_cast_373_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_373_inst_req_1;
      type_cast_373_inst_ack_1<= rack(0);
      type_cast_373_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_373_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext489_525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_373_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_388_inst_req_0;
      type_cast_388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_388_inst_req_1;
      type_cast_388_inst_ack_1<= rack(0);
      type_cast_388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call116_385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv117_389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_401_inst_req_0;
      type_cast_401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_401_inst_req_1;
      type_cast_401_inst_ack_1<= rack(0);
      type_cast_401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call120_398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_419_inst_req_0;
      type_cast_419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_419_inst_req_1;
      type_cast_419_inst_ack_1<= rack(0);
      type_cast_419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call126_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv128_420,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_437_inst_req_0;
      type_cast_437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_437_inst_req_1;
      type_cast_437_inst_ack_1<= rack(0);
      type_cast_437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call132_434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_43_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_43_inst_req_0;
      type_cast_43_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_43_inst_req_1;
      type_cast_43_inst_ack_1<= rack(0);
      type_cast_43_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_43_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_40,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_44,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_455_inst_req_0;
      type_cast_455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_455_inst_req_1;
      type_cast_455_inst_ack_1<= rack(0);
      type_cast_455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call138_452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_473_inst_req_0;
      type_cast_473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_473_inst_req_1;
      type_cast_473_inst_ack_1<= rack(0);
      type_cast_473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call144_470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_491_inst_req_0;
      type_cast_491_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_491_inst_req_1;
      type_cast_491_inst_ack_1<= rack(0);
      type_cast_491_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_491_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call150_488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv152_492,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_509_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_509_inst_req_0;
      type_cast_509_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_509_inst_req_1;
      type_cast_509_inst_ack_1<= rack(0);
      type_cast_509_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_509_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call156_506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_510,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_55_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_55_inst_req_0;
      type_cast_55_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_55_inst_req_1;
      type_cast_55_inst_ack_1<= rack(0);
      type_cast_55_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_55_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_52,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_56,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_567_inst_req_0;
      type_cast_567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_567_inst_req_1;
      type_cast_567_inst_ack_1<= rack(0);
      type_cast_567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp481x_xop_564,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_33_568,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_595_inst_req_0;
      type_cast_595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_595_inst_req_1;
      type_cast_595_inst_ack_1<= rack(0);
      type_cast_595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext477_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_595_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_610_inst_req_0;
      type_cast_610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_610_inst_req_1;
      type_cast_610_inst_ack_1<= rack(0);
      type_cast_610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call172_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_623_inst_req_0;
      type_cast_623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_623_inst_req_1;
      type_cast_623_inst_ack_1<= rack(0);
      type_cast_623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call176_620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv178_624,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_641_inst_req_0;
      type_cast_641_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_641_inst_req_1;
      type_cast_641_inst_ack_1<= rack(0);
      type_cast_641_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_641_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call182_638,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv184_642,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_659_inst_req_0;
      type_cast_659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_659_inst_req_1;
      type_cast_659_inst_ack_1<= rack(0);
      type_cast_659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call188_656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv190_660,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_677_inst_req_0;
      type_cast_677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_677_inst_req_1;
      type_cast_677_inst_ack_1<= rack(0);
      type_cast_677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call194_674,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv196_678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_68_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_68_inst_req_0;
      type_cast_68_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_68_inst_req_1;
      type_cast_68_inst_ack_1<= rack(0);
      type_cast_68_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_68_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_65,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_69,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_695_inst_req_0;
      type_cast_695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_695_inst_req_1;
      type_cast_695_inst_ack_1<= rack(0);
      type_cast_695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call200_692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv202_696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_713_inst_req_0;
      type_cast_713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_713_inst_req_1;
      type_cast_713_inst_ack_1<= rack(0);
      type_cast_713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call206_710,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv208_714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_731_inst_req_0;
      type_cast_731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_731_inst_req_1;
      type_cast_731_inst_ack_1<= rack(0);
      type_cast_731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call212_728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv214_732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_80_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_80_inst_req_0;
      type_cast_80_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_80_inst_req_1;
      type_cast_80_inst_ack_1<= rack(0);
      type_cast_80_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_80_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_77,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_81,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_822_inst_req_0;
      type_cast_822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_822_inst_req_1;
      type_cast_822_inst_ack_1<= rack(0);
      type_cast_822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_822_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2502_1291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_822_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_827_inst_req_0;
      type_cast_827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_827_inst_req_1;
      type_cast_827_inst_ack_1<= rack(0);
      type_cast_827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_827_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x0_980,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_827_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_832_inst_req_0;
      type_cast_832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_832_inst_req_1;
      type_cast_832_inst_ack_1<= rack(0);
      type_cast_832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_832_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x0504_1263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_832_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_837_inst_req_0;
      type_cast_837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_837_inst_req_1;
      type_cast_837_inst_ack_1<= rack(0);
      type_cast_837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_837_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x2_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_837_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_842_inst_req_0;
      type_cast_842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_842_inst_req_1;
      type_cast_842_inst_ack_1<= rack(0);
      type_cast_842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_842_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x2_1343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_842_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_847_inst_req_0;
      type_cast_847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_847_inst_req_1;
      type_cast_847_inst_ack_1<= rack(0);
      type_cast_847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_847_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x1_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv233_848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_870_inst_req_0;
      type_cast_870_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_870_inst_req_1;
      type_cast_870_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen_exec_guard_863(0);
      type_cast_870_inst_gI: SplitGuardInterface generic map(name => "type_cast_870_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_866_delayed_1_0_866,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom240_871,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_893_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_893_inst_req_0;
      type_cast_893_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_893_inst_req_1;
      type_cast_893_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen_exec_guard_863(0);
      type_cast_893_inst_gI: SplitGuardInterface generic map(name => "type_cast_893_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_893_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_893_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_883_delayed_1_0_889,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom244_894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_93_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_93_inst_req_0;
      type_cast_93_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_93_inst_req_1;
      type_cast_93_inst_ack_1<= rack(0);
      type_cast_93_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_93_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_90,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_94,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_953_inst_req_0;
      type_cast_953_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_953_inst_req_1;
      type_cast_953_inst_ack_1<= rack(0);
      type_cast_953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_933_933_delayed_1_0_954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_958_inst
    process(inc251_942) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc251_942(15 downto 0);
      type_cast_958_wire <= tmp_var; -- 
    end process;
    type_cast_968_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_968_inst_req_0;
      type_cast_968_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_968_inst_req_1;
      type_cast_968_inst_ack_1<= rack(0);
      type_cast_968_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_968_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_945_945_delayed_1_0_969,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_973_inst
    process(inc249_932) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc249_932(15 downto 0);
      type_cast_973_wire <= tmp_var; -- 
    end process;
    type_cast_983_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_983_inst_req_0;
      type_cast_983_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_983_inst_req_1;
      type_cast_983_inst_ack_1<= rack(0);
      type_cast_983_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_983_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x1_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_957_957_delayed_1_0_984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_988_inst
    process(inc247_922) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc247_922(15 downto 0);
      type_cast_988_wire <= tmp_var; -- 
    end process;
    type_cast_999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_999_inst_req_0;
      type_cast_999_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_999_inst_req_1;
      type_cast_999_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xend_exec_guard_950(0);
      type_cast_999_inst_gI: SplitGuardInterface generic map(name => "type_cast_999_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_999_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x0_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_1000,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1079_index_1_rename
    process(R_idxprom268_1078_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom268_1078_resized;
      ov(13 downto 0) := iv;
      R_idxprom268_1078_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1079_index_1_resize
    process(idxprom268_1074) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom268_1074;
      ov := iv(13 downto 0);
      R_idxprom268_1078_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1079_root_address_inst
    process(array_obj_ref_1079_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1079_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1079_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1102_index_1_rename
    process(R_idxprom272_1101_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom272_1101_resized;
      ov(13 downto 0) := iv;
      R_idxprom272_1101_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1102_index_1_resize
    process(idxprom272_1097) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom272_1097;
      ov := iv(13 downto 0);
      R_idxprom272_1101_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1102_root_address_inst
    process(array_obj_ref_1102_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1102_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1102_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1538_index_1_rename
    process(R_indvar_1537_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1537_resized;
      ov(13 downto 0) := iv;
      R_indvar_1537_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1538_index_1_resize
    process(indvar_1526) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1526;
      ov := iv(13 downto 0);
      R_indvar_1537_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1538_root_address_inst
    process(array_obj_ref_1538_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1538_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1538_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_380_index_1_rename
    process(R_indvar488_379_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar488_379_resized;
      ov(13 downto 0) := iv;
      R_indvar488_379_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_380_index_1_resize
    process(indvar488_370) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar488_370;
      ov := iv(13 downto 0);
      R_indvar488_379_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_380_root_address_inst
    process(array_obj_ref_380_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_380_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_380_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_602_index_1_rename
    process(R_indvar476_601_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar476_601_resized;
      ov(13 downto 0) := iv;
      R_indvar476_601_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_602_index_1_resize
    process(indvar476_592) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar476_592;
      ov := iv(13 downto 0);
      R_indvar476_601_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_602_root_address_inst
    process(array_obj_ref_602_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_602_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_602_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_rename
    process(R_idxprom240_875_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom240_875_resized;
      ov(13 downto 0) := iv;
      R_idxprom240_875_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_resize
    process(idxprom240_871) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom240_871;
      ov := iv(13 downto 0);
      R_idxprom240_875_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_root_address_inst
    process(array_obj_ref_876_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_876_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_876_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_899_index_1_rename
    process(R_idxprom244_898_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom244_898_resized;
      ov(13 downto 0) := iv;
      R_idxprom244_898_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_899_index_1_resize
    process(idxprom244_894) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom244_894;
      ov := iv(13 downto 0);
      R_idxprom244_898_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_899_root_address_inst
    process(array_obj_ref_899_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_899_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_899_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_addr_0
    process(ptr_deref_1088_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1088_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_base_resize
    process(arrayidx269_1081) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_1081;
      ov := iv(13 downto 0);
      ptr_deref_1088_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_gather_scatter
    process(ptr_deref_1088_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_data_0;
      ov(63 downto 0) := iv;
      tmp270_1089 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_root_address_inst
    process(ptr_deref_1088_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1088_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_addr_0
    process(ptr_deref_1113_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1113_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1113_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_base_resize
    process(arrayidx273_1043_delayed_6_0_1110) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx273_1043_delayed_6_0_1110;
      ov := iv(13 downto 0);
      ptr_deref_1113_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_gather_scatter
    process(tmp270_1089) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp270_1089;
      ov(63 downto 0) := iv;
      ptr_deref_1113_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_root_address_inst
    process(ptr_deref_1113_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1113_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1113_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_addr_0
    process(ptr_deref_1543_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1543_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1543_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_base_resize
    process(arrayidx385_1540) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx385_1540;
      ov := iv(13 downto 0);
      ptr_deref_1543_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_gather_scatter
    process(ptr_deref_1543_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1543_data_0;
      ov(63 downto 0) := iv;
      tmp386_1544 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_root_address_inst
    process(ptr_deref_1543_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1543_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1543_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_517_addr_0
    process(ptr_deref_517_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_517_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_517_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_517_base_resize
    process(arrayidx_382) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_382;
      ov := iv(13 downto 0);
      ptr_deref_517_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_517_gather_scatter
    process(add159_515) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add159_515;
      ov(63 downto 0) := iv;
      ptr_deref_517_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_517_root_address_inst
    process(ptr_deref_517_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_517_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_517_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_739_addr_0
    process(ptr_deref_739_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_739_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_739_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_739_base_resize
    process(arrayidx219_604) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx219_604;
      ov := iv(13 downto 0);
      ptr_deref_739_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_739_gather_scatter
    process(add215_737) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add215_737;
      ov(63 downto 0) := iv;
      ptr_deref_739_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_739_root_address_inst
    process(ptr_deref_739_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_739_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_739_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_addr_0
    process(ptr_deref_885_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_885_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_885_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_base_resize
    process(arrayidx241_878) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx241_878;
      ov := iv(13 downto 0);
      ptr_deref_885_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_gather_scatter
    process(ptr_deref_885_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_885_data_0;
      ov(63 downto 0) := iv;
      tmp242_886 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_root_address_inst
    process(ptr_deref_885_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_885_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_885_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_addr_0
    process(ptr_deref_910_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_910_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_910_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_base_resize
    process(arrayidx245_894_delayed_6_0_907) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx245_894_delayed_6_0_907;
      ov := iv(13 downto 0);
      ptr_deref_910_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_gather_scatter
    process(tmp242_886) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp242_886;
      ov(63 downto 0) := iv;
      ptr_deref_910_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_root_address_inst
    process(ptr_deref_910_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_910_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_910_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_368_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_536_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_368_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_368_branch_req_0,
          ack0 => do_while_stmt_368_branch_ack_0,
          ack1 => do_while_stmt_368_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    do_while_stmt_590_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_758_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_590_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_590_branch_req_0,
          ack0 => do_while_stmt_590_branch_ack_0,
          ack1 => do_while_stmt_590_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    do_while_stmt_817_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1358_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_817_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_817_branch_req_0,
          ack0 => do_while_stmt_817_branch_ack_0,
          ack1 => do_while_stmt_817_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1359_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ifx_xend297_whilex_xend_taken_1355;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1359_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1359_branch_req_0,
          ack0 => if_stmt_1359_branch_ack_0,
          ack1 => if_stmt_1359_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1488_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp378460_1487;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1488_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1488_branch_req_0,
          ack0 => if_stmt_1488_branch_ack_0,
          ack1 => if_stmt_1488_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1654_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1653;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1654_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1654_branch_req_0,
          ack0 => if_stmt_1654_branch_ack_0,
          ack1 => if_stmt_1654_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_298_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp467_297;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_298_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_298_branch_req_0,
          ack0 => if_stmt_298_branch_ack_0,
          ack1 => if_stmt_298_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_313_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp167463_312;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_313_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_313_branch_req_0,
          ack0 => if_stmt_313_branch_ack_0,
          ack1 => if_stmt_313_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_537_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= forx_xbody_forx_xcond163x_xpreheaderx_xloopexit_taken_533;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_537_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_537_branch_req_0,
          ack0 => if_stmt_537_branch_ack_0,
          ack1 => if_stmt_537_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_759_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= forx_xbody169_forx_xend223x_xloopexit_taken_755;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_759_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_759_branch_req_0,
          ack0 => if_stmt_759_branch_ack_0,
          ack1 => if_stmt_759_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1124_inst
    process(count_inp2x_x1_1049_delayed_3_0_1118) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_inp2x_x1_1049_delayed_3_0_1118, type_cast_1123_wire_constant, tmp_var);
      inc275_1125 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1134_inst
    process(add_inp2x_x1_1056_delayed_3_0_1128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp2x_x1_1056_delayed_3_0_1128, type_cast_1133_wire_constant, tmp_var);
      inc277_1135 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1144_inst
    process(add_outx_x0_1063_delayed_2_0_1138) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_outx_x0_1063_delayed_2_0_1138, type_cast_1143_wire_constant, tmp_var);
      inc279_1145 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_921_inst
    process(count_inp1x_x1_900_delayed_1_0_915) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_inp1x_x1_900_delayed_1_0_915, type_cast_920_wire_constant, tmp_var);
      inc247_922 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_931_inst
    process(add_inp1x_x1_907_delayed_1_0_925) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp1x_x1_907_delayed_1_0_925, type_cast_930_wire_constant, tmp_var);
      inc249_932 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_941_inst
    process(add_outx_x1_914_delayed_1_0_935) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_outx_x1_914_delayed_1_0_935, type_cast_940_wire_constant, tmp_var);
      inc251_942 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1505_inst
    process(shr301_787) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr301_787, type_cast_1504_wire_constant, tmp_var);
      tmp471x_xop_1506 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_341_inst
    process(tmp493_330) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp493_330, type_cast_340_wire_constant, tmp_var);
      tmp493x_xop_342 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_563_inst
    process(tmp481_552) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp481_552, type_cast_562_wire_constant, tmp_var);
      tmp481x_xop_564 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1515_inst
    process(iNsTr_81_1510) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_81_1510, type_cast_1514_wire_constant, tmp_var);
      xx_xop_1516 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1647_inst
    process(indvar_1526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1526, type_cast_1646_wire_constant, tmp_var);
      indvarx_xnext_1648 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_351_inst
    process(iNsTr_19_346) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_19_346, type_cast_350_wire_constant, tmp_var);
      xx_xop501_352 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_524_inst
    process(indvar488_370) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar488_370, type_cast_523_wire_constant, tmp_var);
      indvarx_xnext489_525 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_573_inst
    process(iNsTr_33_568) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_33_568, type_cast_572_wire_constant, tmp_var);
      xx_xop500_574 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_746_inst
    process(indvar476_592) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar476_592, type_cast_745_wire_constant, tmp_var);
      indvarx_xnext477_747 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1016_inst
    process(ifx_xend_exec_guard_975_delayed_1_0_1012, cmp257_1009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend_exec_guard_975_delayed_1_0_1012, cmp257_1009, tmp_var);
      ifx_xend_landx_xlhsx_xtrue_taken_1017 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1025_inst
    process(ifx_xend_exec_guard_980_delayed_1_0_1020, NOT_u1_u1_1024_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend_exec_guard_980_delayed_1_0_1020, NOT_u1_u1_1024_wire, tmp_var);
      ifx_xend_ifx_xend297_taken_1026 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1053_inst
    process(landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049, cmp264_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049, cmp264_1046, tmp_var);
      landx_xlhsx_xtrue_ifx_xthen266_taken_1054 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1062_inst
    process(landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057, NOT_u1_u1_1061_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057, NOT_u1_u1_1061_wire, tmp_var);
      landx_xlhsx_xtrue_landx_xlhsx_xtrue288_taken_1063 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1219_inst
    process(landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1215, cmp294_1212) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue288_exec_guard_1124_delayed_1_0_1215, cmp294_1212, tmp_var);
      landx_xlhsx_xtrue288_ifx_xthen296_taken_1220 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1228_inst
    process(landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1223, NOT_u1_u1_1227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue288_exec_guard_1129_delayed_1_0_1223, NOT_u1_u1_1227_wire, tmp_var);
      landx_xlhsx_xtrue288_ifx_xend297_taken_1229 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_274_inst
    process(mul91_264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul91_264, type_cast_273_wire_constant, tmp_var);
      conv102_275 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_285_inst
    process(mul98_269) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul98_269, type_cast_284_wire_constant, tmp_var);
      conv108_286 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1008_inst
    process(conv253_1000, shr236454_775) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv253_1000, shr236454_775, tmp_var);
      cmp257_1009 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1211_inst
    process(conv290_1203, shr263458_781) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv290_1203, shr263458_781, tmp_var);
      cmp294_1212 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1351_inst
    process(conv299_1347, shr301_787) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv299_1347, shr301_787, tmp_var);
      cmp302_1352 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1652_inst
    process(indvarx_xnext_1648, tmp475_1523) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1648, tmp475_1523, tmp_var);
      exitcond1_1653 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_529_inst
    process(indvarx_xnext489_525, tmp498_359) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext489_525, tmp498_359, tmp_var);
      exitcond2_530 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_751_inst
    process(indvarx_xnext477_747, tmp486_581) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext477_747, tmp486_581, tmp_var);
      exitcond_752 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_329_inst
    process(tmp492_324) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp492_324, type_cast_328_wire_constant, tmp_var);
      tmp493_330 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_551_inst
    process(tmp480_546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp480_546, type_cast_550_wire_constant, tmp_var);
      tmp481_552 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_774_inst
    process(conv102_275) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv102_275, type_cast_773_wire_constant, tmp_var);
      shr236454_775 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_780_inst
    process(conv108_286) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv108_286, type_cast_779_wire_constant, tmp_var);
      shr263458_781 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_786_inst
    process(mul85_259) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul85_259, type_cast_785_wire_constant, tmp_var);
      shr301_787 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1391_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1390_wire_constant, tmp_var);
      shr317_1392 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1401_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1400_wire_constant, tmp_var);
      shr323_1402 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1411_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1410_wire_constant, tmp_var);
      shr329_1412 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1421_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1420_wire_constant, tmp_var);
      shr335_1422 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1431_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1430_wire_constant, tmp_var);
      shr341_1432 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1441_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1440_wire_constant, tmp_var);
      shr347_1442 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1451_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1450_wire_constant, tmp_var);
      shr353_1452 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1553_inst
    process(tmp386_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp386_1544, type_cast_1552_wire_constant, tmp_var);
      shr393_1554 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1563_inst
    process(tmp386_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp386_1544, type_cast_1562_wire_constant, tmp_var);
      shr399_1564 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1573_inst
    process(tmp386_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp386_1544, type_cast_1572_wire_constant, tmp_var);
      shr405_1574 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1583_inst
    process(tmp386_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp386_1544, type_cast_1582_wire_constant, tmp_var);
      shr411_1584 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1593_inst
    process(tmp386_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp386_1544, type_cast_1592_wire_constant, tmp_var);
      shr417_1594 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1603_inst
    process(tmp386_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp386_1544, type_cast_1602_wire_constant, tmp_var);
      shr423_1604 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1613_inst
    process(tmp386_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp386_1544, type_cast_1612_wire_constant, tmp_var);
      shr429_1614 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_253_inst
    process(add66_224, add57_199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add66_224, add57_199, tmp_var);
      mul_254 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_258_inst
    process(mul_254, add75_249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_254, add75_249, tmp_var);
      mul85_259 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_263_inst
    process(add21_99, add12_74) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add21_99, add12_74, tmp_var);
      mul91_264 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_268_inst
    process(add48_174, add39_149) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add48_174, add39_149, tmp_var);
      mul98_269 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_279_inst
    process(conv102_275, add_49) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv102_275, add_49, tmp_var);
      mul105_280 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_290_inst
    process(conv108_286, add30_124) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv108_286, add30_124, tmp_var);
      mul111_291 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_323_inst
    process(add_49, conv102_275) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_49, conv102_275, tmp_var);
      tmp492_324 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_545_inst
    process(add30_124, conv108_286) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add30_124, conv108_286, tmp_var);
      tmp480_546 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1024_inst
    process(cmp257_1009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp257_1009, tmp_var);
      NOT_u1_u1_1024_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1061_inst
    process(cmp264_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp264_1046, tmp_var);
      NOT_u1_u1_1061_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1227_inst
    process(cmp294_1212) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp294_1212, tmp_var);
      NOT_u1_u1_1227_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1358_inst
    process(cmp302_1352) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp302_1352, tmp_var);
      NOT_u1_u1_1358_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_536_inst
    process(exitcond2_530) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", exitcond2_530, tmp_var);
      NOT_u1_u1_536_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_758_inst
    process(exitcond_752) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", exitcond_752, tmp_var);
      NOT_u1_u1_758_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_859_inst
    process(cmp237_853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp237_853, tmp_var);
      whilex_xbody_ifx_xend_taken_860 <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1152_inst
    process(ifx_xthen266_landx_xlhsx_xtrue288_taken_1148, landx_xlhsx_xtrue_landx_xlhsx_xtrue288_taken_1063) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xthen266_landx_xlhsx_xtrue288_taken_1148, landx_xlhsx_xtrue_landx_xlhsx_xtrue288_taken_1063, tmp_var);
      landx_xlhsx_xtrue288_exec_guard_1153 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_949_inst
    process(ifx_xthen_ifx_xend_taken_945, whilex_xbody_ifx_xend_taken_860) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xthen_ifx_xend_taken_945, whilex_xbody_ifx_xend_taken_860, tmp_var);
      ifx_xend_exec_guard_950 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_123_inst
    process(shl27_112, conv29_119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_112, conv29_119, tmp_var);
      add30_124 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_148_inst
    process(shl36_137, conv38_144) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_137, conv38_144, tmp_var);
      add39_149 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_173_inst
    process(shl45_162, conv47_169) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_162, conv47_169, tmp_var);
      add48_174 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_198_inst
    process(shl54_187, conv56_194) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_187, conv56_194, tmp_var);
      add57_199 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_223_inst
    process(shl63_212, conv65_219) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl63_212, conv65_219, tmp_var);
      add66_224 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_248_inst
    process(shl72_237, conv74_244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl72_237, conv74_244, tmp_var);
      add75_249 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_48_inst
    process(shl_37, conv3_44) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_37, conv3_44, tmp_var);
      add_49 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_73_inst
    process(shl9_62, conv11_69) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_62, conv11_69, tmp_var);
      add12_74 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_98_inst
    process(shl18_87, conv20_94) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_87, conv20_94, tmp_var);
      add21_99 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_406_inst
    process(shl119_395, conv122_402) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl119_395, conv122_402, tmp_var);
      add123_407 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_424_inst
    process(shl125_413, conv128_420) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl125_413, conv128_420, tmp_var);
      add129_425 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_442_inst
    process(shl131_431, conv134_438) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl131_431, conv134_438, tmp_var);
      add135_443 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_460_inst
    process(shl137_449, conv140_456) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl137_449, conv140_456, tmp_var);
      add141_461 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_478_inst
    process(shl143_467, conv146_474) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl143_467, conv146_474, tmp_var);
      add147_479 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_496_inst
    process(shl149_485, conv152_492) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl149_485, conv152_492, tmp_var);
      add153_497 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_514_inst
    process(shl155_503, conv158_510) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl155_503, conv158_510, tmp_var);
      add159_515 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_628_inst
    process(shl175_617, conv178_624) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl175_617, conv178_624, tmp_var);
      add179_629 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_646_inst
    process(shl181_635, conv184_642) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl181_635, conv184_642, tmp_var);
      add185_647 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_664_inst
    process(shl187_653, conv190_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl187_653, conv190_660, tmp_var);
      add191_665 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_682_inst
    process(shl193_671, conv196_678) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl193_671, conv196_678, tmp_var);
      add197_683 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_700_inst
    process(shl199_689, conv202_696) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl199_689, conv202_696, tmp_var);
      add203_701 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_718_inst
    process(shl205_707, conv208_714) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl205_707, conv208_714, tmp_var);
      add209_719 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_736_inst
    process(shl211_725, conv214_732) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl211_725, conv214_732, tmp_var);
      add215_737 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_111_inst
    process(conv26_106) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_106, type_cast_110_wire_constant, tmp_var);
      shl27_112 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_136_inst
    process(conv35_131) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_131, type_cast_135_wire_constant, tmp_var);
      shl36_137 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_161_inst
    process(conv44_156) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_156, type_cast_160_wire_constant, tmp_var);
      shl45_162 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_186_inst
    process(conv53_181) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_181, type_cast_185_wire_constant, tmp_var);
      shl54_187 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_211_inst
    process(conv62_206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv62_206, type_cast_210_wire_constant, tmp_var);
      shl63_212 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_236_inst
    process(conv71_231) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv71_231, type_cast_235_wire_constant, tmp_var);
      shl72_237 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_36_inst
    process(conv1_31) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_31, type_cast_35_wire_constant, tmp_var);
      shl_37 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_61_inst
    process(conv8_56) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_56, type_cast_60_wire_constant, tmp_var);
      shl9_62 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_86_inst
    process(conv17_81) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_81, type_cast_85_wire_constant, tmp_var);
      shl18_87 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_394_inst
    process(conv117_389) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv117_389, type_cast_393_wire_constant, tmp_var);
      shl119_395 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_412_inst
    process(add123_407) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add123_407, type_cast_411_wire_constant, tmp_var);
      shl125_413 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_430_inst
    process(add129_425) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add129_425, type_cast_429_wire_constant, tmp_var);
      shl131_431 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_448_inst
    process(add135_443) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add135_443, type_cast_447_wire_constant, tmp_var);
      shl137_449 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_466_inst
    process(add141_461) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add141_461, type_cast_465_wire_constant, tmp_var);
      shl143_467 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_484_inst
    process(add147_479) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add147_479, type_cast_483_wire_constant, tmp_var);
      shl149_485 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_502_inst
    process(add153_497) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add153_497, type_cast_501_wire_constant, tmp_var);
      shl155_503 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_616_inst
    process(conv173_611) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv173_611, type_cast_615_wire_constant, tmp_var);
      shl175_617 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_634_inst
    process(add179_629) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add179_629, type_cast_633_wire_constant, tmp_var);
      shl181_635 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_652_inst
    process(add185_647) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add185_647, type_cast_651_wire_constant, tmp_var);
      shl187_653 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_670_inst
    process(add191_665) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add191_665, type_cast_669_wire_constant, tmp_var);
      shl193_671 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_688_inst
    process(add197_683) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add197_683, type_cast_687_wire_constant, tmp_var);
      shl199_689 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_706_inst
    process(add203_701) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add203_701, type_cast_705_wire_constant, tmp_var);
      shl205_707 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_724_inst
    process(add209_719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add209_719, type_cast_723_wire_constant, tmp_var);
      shl211_725 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1381_inst
    process(conv308_1377, conv226_1369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv308_1377, conv226_1369, tmp_var);
      sub_1382 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1486_inst
    process(mul85_259) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul85_259, type_cast_1485_wire_constant, tmp_var);
      cmp378460_1487 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1499_inst
    process(shr301_787) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr301_787, type_cast_1498_wire_constant, tmp_var);
      tmp472_1500 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_296_inst
    process(mul105_280) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul105_280, type_cast_295_wire_constant, tmp_var);
      cmp467_297 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_311_inst
    process(mul111_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul111_291, type_cast_310_wire_constant, tmp_var);
      cmp167463_312 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_335_inst
    process(tmp493_330) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp493_330, type_cast_334_wire_constant, tmp_var);
      tmp494_336 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_557_inst
    process(tmp481_552) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp481_552, type_cast_556_wire_constant, tmp_var);
      tmp482_558 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1045_inst
    process(conv260_1037, shr263458_781) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv260_1037, shr263458_781, tmp_var);
      cmp264_1046 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_852_inst
    process(conv233_848, shr236454_775) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv233_848, shr236454_775, tmp_var);
      cmp237_853 <= tmp_var; --
    end process;
    -- shared split operator group (120) : array_obj_ref_1079_index_offset 
    ApIntAdd_group_120: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom268_1078_scaled;
      array_obj_ref_1079_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1079_index_offset_req_0;
      array_obj_ref_1079_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1079_index_offset_req_1;
      array_obj_ref_1079_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_120_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_120_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_120",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 120
    -- shared split operator group (121) : array_obj_ref_1102_index_offset 
    ApIntAdd_group_121: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom272_1101_scaled;
      array_obj_ref_1102_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1102_index_offset_req_0;
      array_obj_ref_1102_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1102_index_offset_req_1;
      array_obj_ref_1102_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_121_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_121_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_121",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 121
    -- shared split operator group (122) : array_obj_ref_1538_index_offset 
    ApIntAdd_group_122: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1537_scaled;
      array_obj_ref_1538_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1538_index_offset_req_0;
      array_obj_ref_1538_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1538_index_offset_req_1;
      array_obj_ref_1538_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_122_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_122_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : array_obj_ref_380_index_offset 
    ApIntAdd_group_123: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar488_379_scaled;
      array_obj_ref_380_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_380_index_offset_req_0;
      array_obj_ref_380_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_380_index_offset_req_1;
      array_obj_ref_380_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_123_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_123_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : array_obj_ref_602_index_offset 
    ApIntAdd_group_124: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar476_601_scaled;
      array_obj_ref_602_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_602_index_offset_req_0;
      array_obj_ref_602_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_602_index_offset_req_1;
      array_obj_ref_602_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_124_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_124_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : array_obj_ref_876_index_offset 
    ApIntAdd_group_125: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom240_875_scaled;
      array_obj_ref_876_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_876_index_offset_req_0;
      array_obj_ref_876_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_876_index_offset_req_1;
      array_obj_ref_876_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_125_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_125_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- shared split operator group (126) : array_obj_ref_899_index_offset 
    ApIntAdd_group_126: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom244_898_scaled;
      array_obj_ref_899_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_899_index_offset_req_0;
      array_obj_ref_899_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_899_index_offset_req_1;
      array_obj_ref_899_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_126_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_126_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_126",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 126
    -- unary operator type_cast_1367_inst
    process(call225_768) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call225_768, tmp_var);
      type_cast_1367_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1375_inst
    process(call307_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call307_1372, tmp_var);
      type_cast_1375_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1088_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1088_load_0_req_0;
      ptr_deref_1088_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1088_load_0_req_1;
      ptr_deref_1088_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xthen266_exec_guard_1025_delayed_7_0_1084(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1088_word_address_0;
      ptr_deref_1088_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1543_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1543_load_0_req_0;
      ptr_deref_1543_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1543_load_0_req_1;
      ptr_deref_1543_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1543_word_address_0;
      ptr_deref_1543_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_885_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_885_load_0_req_0;
      ptr_deref_885_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_885_load_0_req_1;
      ptr_deref_885_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xthen_exec_guard_876_delayed_7_0_881(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_885_word_address_0;
      ptr_deref_885_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : ptr_deref_910_store_0 ptr_deref_1113_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_910_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1113_store_0_req_0;
      ptr_deref_910_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1113_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_910_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1113_store_0_req_1;
      ptr_deref_910_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1113_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xthen266_exec_guard_1042_delayed_13_0_1107(0);
      guard_vector(1)  <= ifx_xthen_exec_guard_893_delayed_13_0_904(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_910_word_address_0 & ptr_deref_1113_word_address_0;
      data_in <= ptr_deref_910_data_0 & ptr_deref_1113_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_517_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_517_store_0_req_0;
      ptr_deref_517_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_517_store_0_req_1;
      ptr_deref_517_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_517_word_address_0;
      data_in <= ptr_deref_517_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_739_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_739_store_0_req_0;
      ptr_deref_739_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_739_store_0_req_1;
      ptr_deref_739_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_739_word_address_0;
      data_in <= ptr_deref_739_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Concat_input_pipe_25_inst RPIPE_Concat_input_pipe_39_inst RPIPE_Concat_input_pipe_51_inst RPIPE_Concat_input_pipe_64_inst RPIPE_Concat_input_pipe_76_inst RPIPE_Concat_input_pipe_89_inst RPIPE_Concat_input_pipe_101_inst RPIPE_Concat_input_pipe_114_inst RPIPE_Concat_input_pipe_126_inst RPIPE_Concat_input_pipe_139_inst RPIPE_Concat_input_pipe_151_inst RPIPE_Concat_input_pipe_164_inst RPIPE_Concat_input_pipe_176_inst RPIPE_Concat_input_pipe_189_inst RPIPE_Concat_input_pipe_201_inst RPIPE_Concat_input_pipe_214_inst RPIPE_Concat_input_pipe_226_inst RPIPE_Concat_input_pipe_239_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(143 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 17 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 17 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 17 downto 0);
      signal guard_vector : std_logic_vector( 17 downto 0);
      constant outBUFs : IntegerArray(17 downto 0) := (17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(17 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false);
      constant guardBuffering: IntegerArray(17 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2);
      -- 
    begin -- 
      reqL_unguarded(17) <= RPIPE_Concat_input_pipe_25_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Concat_input_pipe_39_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Concat_input_pipe_51_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Concat_input_pipe_64_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Concat_input_pipe_76_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Concat_input_pipe_89_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Concat_input_pipe_101_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Concat_input_pipe_114_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Concat_input_pipe_126_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Concat_input_pipe_139_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Concat_input_pipe_151_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Concat_input_pipe_164_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Concat_input_pipe_176_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Concat_input_pipe_189_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Concat_input_pipe_201_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Concat_input_pipe_214_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Concat_input_pipe_226_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Concat_input_pipe_239_inst_req_0;
      RPIPE_Concat_input_pipe_25_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Concat_input_pipe_39_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Concat_input_pipe_51_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Concat_input_pipe_64_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Concat_input_pipe_76_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Concat_input_pipe_89_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Concat_input_pipe_101_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Concat_input_pipe_114_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Concat_input_pipe_126_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Concat_input_pipe_139_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Concat_input_pipe_151_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Concat_input_pipe_164_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Concat_input_pipe_176_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Concat_input_pipe_189_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Concat_input_pipe_201_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Concat_input_pipe_214_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Concat_input_pipe_226_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Concat_input_pipe_239_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(17) <= RPIPE_Concat_input_pipe_25_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Concat_input_pipe_39_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Concat_input_pipe_51_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Concat_input_pipe_64_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Concat_input_pipe_76_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Concat_input_pipe_89_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Concat_input_pipe_101_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Concat_input_pipe_114_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Concat_input_pipe_126_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Concat_input_pipe_139_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Concat_input_pipe_151_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Concat_input_pipe_164_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Concat_input_pipe_176_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Concat_input_pipe_189_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Concat_input_pipe_201_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Concat_input_pipe_214_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Concat_input_pipe_226_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Concat_input_pipe_239_inst_req_1;
      RPIPE_Concat_input_pipe_25_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Concat_input_pipe_39_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Concat_input_pipe_51_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Concat_input_pipe_64_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Concat_input_pipe_76_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Concat_input_pipe_89_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Concat_input_pipe_101_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Concat_input_pipe_114_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Concat_input_pipe_126_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Concat_input_pipe_139_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Concat_input_pipe_151_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Concat_input_pipe_164_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Concat_input_pipe_176_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Concat_input_pipe_189_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Concat_input_pipe_201_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Concat_input_pipe_214_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Concat_input_pipe_226_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Concat_input_pipe_239_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      call_26 <= data_out(143 downto 136);
      call2_40 <= data_out(135 downto 128);
      call5_52 <= data_out(127 downto 120);
      call10_65 <= data_out(119 downto 112);
      call14_77 <= data_out(111 downto 104);
      call19_90 <= data_out(103 downto 96);
      call23_102 <= data_out(95 downto 88);
      call28_115 <= data_out(87 downto 80);
      call32_127 <= data_out(79 downto 72);
      call37_140 <= data_out(71 downto 64);
      call41_152 <= data_out(63 downto 56);
      call46_165 <= data_out(55 downto 48);
      call50_177 <= data_out(47 downto 40);
      call55_190 <= data_out(39 downto 32);
      call59_202 <= data_out(31 downto 24);
      call64_215 <= data_out(23 downto 16);
      call68_227 <= data_out(15 downto 8);
      call73_240 <= data_out(7 downto 0);
      Concat_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "Concat_input_pipe_read_0_gI", nreqs => 18, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Concat_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "Concat_input_pipe_read_0", data_width => 8,  num_reqs => 18,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Concat_input_pipe_pipe_read_req(1),
          oack => Concat_input_pipe_pipe_read_ack(1),
          odata => Concat_input_pipe_pipe_read_data(15 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Concat_input_pipe_384_inst RPIPE_Concat_input_pipe_397_inst RPIPE_Concat_input_pipe_415_inst RPIPE_Concat_input_pipe_433_inst RPIPE_Concat_input_pipe_451_inst RPIPE_Concat_input_pipe_469_inst RPIPE_Concat_input_pipe_487_inst RPIPE_Concat_input_pipe_505_inst RPIPE_Concat_input_pipe_606_inst RPIPE_Concat_input_pipe_619_inst RPIPE_Concat_input_pipe_637_inst RPIPE_Concat_input_pipe_655_inst RPIPE_Concat_input_pipe_673_inst RPIPE_Concat_input_pipe_691_inst RPIPE_Concat_input_pipe_709_inst RPIPE_Concat_input_pipe_727_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 15 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= RPIPE_Concat_input_pipe_384_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Concat_input_pipe_397_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Concat_input_pipe_415_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Concat_input_pipe_433_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Concat_input_pipe_451_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Concat_input_pipe_469_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Concat_input_pipe_487_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Concat_input_pipe_505_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Concat_input_pipe_606_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Concat_input_pipe_619_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Concat_input_pipe_637_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Concat_input_pipe_655_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Concat_input_pipe_673_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Concat_input_pipe_691_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Concat_input_pipe_709_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Concat_input_pipe_727_inst_req_0;
      RPIPE_Concat_input_pipe_384_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Concat_input_pipe_397_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Concat_input_pipe_415_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Concat_input_pipe_433_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Concat_input_pipe_451_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Concat_input_pipe_469_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Concat_input_pipe_487_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Concat_input_pipe_505_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Concat_input_pipe_606_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Concat_input_pipe_619_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Concat_input_pipe_637_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Concat_input_pipe_655_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Concat_input_pipe_673_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Concat_input_pipe_691_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Concat_input_pipe_709_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Concat_input_pipe_727_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= RPIPE_Concat_input_pipe_384_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Concat_input_pipe_397_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Concat_input_pipe_415_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Concat_input_pipe_433_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Concat_input_pipe_451_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Concat_input_pipe_469_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Concat_input_pipe_487_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Concat_input_pipe_505_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Concat_input_pipe_606_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Concat_input_pipe_619_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Concat_input_pipe_637_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Concat_input_pipe_655_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Concat_input_pipe_673_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Concat_input_pipe_691_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Concat_input_pipe_709_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Concat_input_pipe_727_inst_req_1;
      RPIPE_Concat_input_pipe_384_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Concat_input_pipe_397_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Concat_input_pipe_415_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Concat_input_pipe_433_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Concat_input_pipe_451_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Concat_input_pipe_469_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Concat_input_pipe_487_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Concat_input_pipe_505_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Concat_input_pipe_606_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Concat_input_pipe_619_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Concat_input_pipe_637_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Concat_input_pipe_655_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Concat_input_pipe_673_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Concat_input_pipe_691_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Concat_input_pipe_709_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Concat_input_pipe_727_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      call116_385 <= data_out(127 downto 120);
      call120_398 <= data_out(119 downto 112);
      call126_416 <= data_out(111 downto 104);
      call132_434 <= data_out(103 downto 96);
      call138_452 <= data_out(95 downto 88);
      call144_470 <= data_out(87 downto 80);
      call150_488 <= data_out(79 downto 72);
      call156_506 <= data_out(71 downto 64);
      call172_607 <= data_out(63 downto 56);
      call176_620 <= data_out(55 downto 48);
      call182_638 <= data_out(47 downto 40);
      call188_656 <= data_out(39 downto 32);
      call194_674 <= data_out(31 downto 24);
      call200_692 <= data_out(23 downto 16);
      call206_710 <= data_out(15 downto 8);
      call212_728 <= data_out(7 downto 0);
      Concat_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "Concat_input_pipe_read_1_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Concat_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "Concat_input_pipe_read_1", data_width => 8,  num_reqs => 16,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Concat_input_pipe_pipe_read_req(0),
          oack => Concat_input_pipe_pipe_read_ack(0),
          odata => Concat_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_Concat_output_pipe_1457_inst WPIPE_Concat_output_pipe_1460_inst WPIPE_Concat_output_pipe_1463_inst WPIPE_Concat_output_pipe_1466_inst WPIPE_Concat_output_pipe_1469_inst WPIPE_Concat_output_pipe_1472_inst WPIPE_Concat_output_pipe_1475_inst WPIPE_Concat_output_pipe_1478_inst WPIPE_Concat_output_pipe_1619_inst WPIPE_Concat_output_pipe_1622_inst WPIPE_Concat_output_pipe_1625_inst WPIPE_Concat_output_pipe_1628_inst WPIPE_Concat_output_pipe_1631_inst WPIPE_Concat_output_pipe_1634_inst WPIPE_Concat_output_pipe_1637_inst WPIPE_Concat_output_pipe_1640_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_Concat_output_pipe_1457_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Concat_output_pipe_1460_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Concat_output_pipe_1463_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Concat_output_pipe_1466_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Concat_output_pipe_1469_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Concat_output_pipe_1472_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Concat_output_pipe_1475_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Concat_output_pipe_1478_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Concat_output_pipe_1619_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Concat_output_pipe_1622_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Concat_output_pipe_1625_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Concat_output_pipe_1628_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Concat_output_pipe_1631_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Concat_output_pipe_1634_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Concat_output_pipe_1637_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Concat_output_pipe_1640_inst_req_0;
      WPIPE_Concat_output_pipe_1457_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1460_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1463_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1466_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1469_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1472_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1475_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1478_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1619_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1622_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1625_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1628_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1631_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1634_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1637_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1640_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_Concat_output_pipe_1457_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Concat_output_pipe_1460_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Concat_output_pipe_1463_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Concat_output_pipe_1466_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Concat_output_pipe_1469_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Concat_output_pipe_1472_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Concat_output_pipe_1475_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Concat_output_pipe_1478_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Concat_output_pipe_1619_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Concat_output_pipe_1622_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Concat_output_pipe_1625_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Concat_output_pipe_1628_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Concat_output_pipe_1631_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Concat_output_pipe_1634_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Concat_output_pipe_1637_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Concat_output_pipe_1640_inst_req_1;
      WPIPE_Concat_output_pipe_1457_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1460_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1463_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1466_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1469_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1472_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1475_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1478_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1619_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1622_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1625_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1628_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1631_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1634_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1637_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1640_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv356_1456 & conv350_1446 & conv344_1436 & conv338_1426 & conv332_1416 & conv326_1406 & conv320_1396 & conv314_1386 & conv432_1618 & conv426_1608 & conv420_1598 & conv414_1588 & conv408_1578 & conv402_1568 & conv396_1558 & conv390_1548;
      Concat_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "Concat_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Concat_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "Concat_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Concat_output_pipe_pipe_write_req(0),
          oack => Concat_output_pipe_pipe_write_ack(0),
          odata => Concat_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_768_call call_stmt_1372_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_768_call_req_0;
      reqL_unguarded(0) <= call_stmt_1372_call_req_0;
      call_stmt_768_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1372_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_768_call_req_1;
      reqR_unguarded(0) <= call_stmt_1372_call_req_1;
      call_stmt_768_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1372_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call225_768 <= data_out(127 downto 64);
      call307_1372 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end concat_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_14_inst_req_0 : boolean;
  signal WPIPE_timer_req_14_inst_ack_0 : boolean;
  signal WPIPE_timer_req_14_inst_req_1 : boolean;
  signal WPIPE_timer_req_14_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_19_inst_req_0 : boolean;
  signal RPIPE_timer_resp_19_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_19_inst_req_1 : boolean;
  signal RPIPE_timer_resp_19_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_sample_start_
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/req
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_sample_start_
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_19_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_14_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_sample_completed_
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_update_start_
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/ack
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/$entry
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_14_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_14_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_update_completed_
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/$exit
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_14_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_update_start_
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_sample_completed_
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/ra
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/$entry
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_19_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_19_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_update_completed_
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/$exit
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_19_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_17_to_assign_stmt_20/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(2) & timer_CP_0_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_16_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_16_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_19_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_19_inst_req_0;
      RPIPE_timer_resp_19_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_19_inst_req_1;
      RPIPE_timer_resp_19_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_14_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_14_inst_req_0;
      WPIPE_timer_req_14_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_14_inst_req_1;
      WPIPE_timer_req_14_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_16_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_3831_start: Boolean;
  signal timerDaemon_CP_3831_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1679_req_1 : boolean;
  signal nCOUNTER_1692_1683_buf_req_0 : boolean;
  signal nCOUNTER_1692_1683_buf_req_1 : boolean;
  signal nCOUNTER_1692_1683_buf_ack_1 : boolean;
  signal RPIPE_timer_req_1686_inst_req_1 : boolean;
  signal RPIPE_timer_req_1686_inst_ack_0 : boolean;
  signal nCOUNTER_1692_1683_buf_ack_0 : boolean;
  signal RPIPE_timer_req_1686_inst_req_0 : boolean;
  signal WPIPE_timer_resp_1694_inst_req_0 : boolean;
  signal RPIPE_timer_req_1686_inst_ack_1 : boolean;
  signal phi_stmt_1679_req_0 : boolean;
  signal do_while_stmt_1677_branch_ack_0 : boolean;
  signal phi_stmt_1679_ack_0 : boolean;
  signal WPIPE_timer_resp_1694_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_1694_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_1694_inst_req_1 : boolean;
  signal do_while_stmt_1677_branch_req_0 : boolean;
  signal do_while_stmt_1677_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_3831_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3831_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_3831_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3831_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_3831: Block -- control-path 
    signal timerDaemon_CP_3831_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_3831_elements(0) <= timerDaemon_CP_3831_start;
    timerDaemon_CP_3831_symbol <= timerDaemon_CP_3831_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1676/$entry
      -- CP-element group 0: 	 branch_block_stmt_1676/do_while_stmt_1677__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1676/branch_block_stmt_1676__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1676/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1676/do_while_stmt_1677__exit__
      -- CP-element group 1: 	 branch_block_stmt_1676/branch_block_stmt_1676__exit__
      -- 
    timerDaemon_CP_3831_elements(1) <= timerDaemon_CP_3831_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1676/do_while_stmt_1677/$entry
      -- CP-element group 2: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677__entry__
      -- 
    timerDaemon_CP_3831_elements(2) <= timerDaemon_CP_3831_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677__exit__
      -- 
    -- Element group timerDaemon_CP_3831_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_back
      -- 
    -- Element group timerDaemon_CP_3831_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1676/do_while_stmt_1677/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_taken/$entry
      -- 
    timerDaemon_CP_3831_elements(5) <= timerDaemon_CP_3831_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_body_done
      -- 
    timerDaemon_CP_3831_elements(6) <= timerDaemon_CP_3831_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_3831_elements(7) <= timerDaemon_CP_3831_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_3831_elements(8) <= timerDaemon_CP_3831_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/loop_body_start
      -- 
    -- Element group timerDaemon_CP_3831_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/condition_evaluated
      -- 
    condition_evaluated_3855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(10), ack => do_while_stmt_1677_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(14) & timerDaemon_CP_3831_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_sample_req
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(9) & timerDaemon_CP_3831_elements(15) & timerDaemon_CP_3831_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_sample_ack
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(17) & timerDaemon_CP_3831_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(16) & timerDaemon_CP_3831_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(18) & timerDaemon_CP_3831_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(9) & timerDaemon_CP_3831_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(9) & timerDaemon_CP_3831_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_3831_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_3831_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_loopback_trigger
      -- 
    timerDaemon_CP_3831_elements(19) <= timerDaemon_CP_3831_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_loopback_sample_req_ps
      -- 
    phi_stmt_1679_loopback_sample_req_3870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1679_loopback_sample_req_3870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(20), ack => phi_stmt_1679_req_1); -- 
    -- Element group timerDaemon_CP_3831_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_entry_trigger
      -- 
    timerDaemon_CP_3831_elements(21) <= timerDaemon_CP_3831_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_entry_sample_req_ps
      -- 
    phi_stmt_1679_entry_sample_req_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1679_entry_sample_req_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(22), ack => phi_stmt_1679_req_0); -- 
    -- Element group timerDaemon_CP_3831_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_phi_mux_ack_ps
      -- 
    phi_stmt_1679_phi_mux_ack_3876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1679_ack_0, ack => timerDaemon_CP_3831_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_3831_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_start__ps
      -- 
    -- Element group timerDaemon_CP_3831_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_completed__ps
      -- 
    timerDaemon_CP_3831_elements(26) <= timerDaemon_CP_3831_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_completed_
      -- 
    -- Element group timerDaemon_CP_3831_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_3831_elements(25), ack => timerDaemon_CP_3831_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_start_
      -- 
    req_3897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(28), ack => nCOUNTER_1692_1683_buf_req_0); -- 
    -- Element group timerDaemon_CP_3831_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_start_
      -- 
    req_3902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(29), ack => nCOUNTER_1692_1683_buf_req_1); -- 
    -- Element group timerDaemon_CP_3831_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_completed_
      -- 
    ack_3898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1692_1683_buf_ack_0, ack => timerDaemon_CP_3831_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_completed__ps
      -- 
    ack_3903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1692_1683_buf_ack_1, ack => timerDaemon_CP_3831_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(9) & timerDaemon_CP_3831_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/$entry
      -- 
    rr_3916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(33), ack => RPIPE_timer_req_1686_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(11) & timerDaemon_CP_3831_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/$entry
      -- 
    cr_3921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(34), ack => RPIPE_timer_req_1686_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(13) & timerDaemon_CP_3831_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/$exit
      -- 
    ra_3917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1686_inst_ack_0, ack => timerDaemon_CP_3831_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/$exit
      -- 
    ca_3922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1686_inst_ack_1, ack => timerDaemon_CP_3831_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/req
      -- 
    req_3930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(37), ack => WPIPE_timer_resp_1694_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(18) & timerDaemon_CP_3831_elements(36) & timerDaemon_CP_3831_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/req
      -- 
    ack_3931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1694_inst_ack_0, ack => timerDaemon_CP_3831_elements(38)); -- 
    req_3935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3831_elements(38), ack => WPIPE_timer_resp_1694_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/ack
      -- 
    ack_3936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1694_inst_ack_1, ack => timerDaemon_CP_3831_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_3831_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_3831_elements(9), ack => timerDaemon_CP_3831_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3831_elements(12) & timerDaemon_CP_3831_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3831_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_exit/ack
      -- 
    ack_3941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1677_branch_ack_0, ack => timerDaemon_CP_3831_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_taken/ack
      -- 
    ack_3945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1677_branch_ack_1, ack => timerDaemon_CP_3831_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1676/do_while_stmt_1677/$exit
      -- 
    timerDaemon_CP_3831_elements(44) <= timerDaemon_CP_3831_elements(3);
    timerDaemon_do_while_stmt_1677_terminator_3946: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1677_terminator_3946", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_3831_elements(6),loop_continue => timerDaemon_CP_3831_elements(43),loop_terminate => timerDaemon_CP_3831_elements(42),loop_back => timerDaemon_CP_3831_elements(4),loop_exit => timerDaemon_CP_3831_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1679_phi_seq_3904_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_3831_elements(21);
      timerDaemon_CP_3831_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_3831_elements(24);
      timerDaemon_CP_3831_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_3831_elements(26);
      timerDaemon_CP_3831_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_3831_elements(19);
      timerDaemon_CP_3831_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_3831_elements(30);
      timerDaemon_CP_3831_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_3831_elements(31);
      timerDaemon_CP_3831_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1679_phi_seq_3904 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1679_phi_seq_3904") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_3831_elements(11), 
          phi_sample_ack => timerDaemon_CP_3831_elements(17), 
          phi_update_req => timerDaemon_CP_3831_elements(13), 
          phi_update_ack => timerDaemon_CP_3831_elements(18), 
          phi_mux_ack => timerDaemon_CP_3831_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3856_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_3831_elements(7);
        preds(1)  <= timerDaemon_CP_3831_elements(8);
        entry_tmerge_3856 : transition_merge -- 
          generic map(name => " entry_tmerge_3856")
          port map (preds => preds, symbol_out => timerDaemon_CP_3831_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1679 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1686_wire : std_logic_vector(0 downto 0);
    signal konst_1690_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1698_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1692 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1692_1683_buffered : std_logic_vector(63 downto 0);
    signal req_1684 : std_logic_vector(0 downto 0);
    signal type_cast_1682_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1690_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1698_wire_constant <= "1";
    type_cast_1682_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1679: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1682_wire_constant & nCOUNTER_1692_1683_buffered;
      req <= phi_stmt_1679_req_0 & phi_stmt_1679_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1679",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1679_ack_0,
          idata => idata,
          odata => COUNTER_1679,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1679
    nCOUNTER_1692_1683_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1692_1683_buf_req_0;
      nCOUNTER_1692_1683_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1692_1683_buf_req_1;
      nCOUNTER_1692_1683_buf_ack_1<= rack(0);
      nCOUNTER_1692_1683_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1692_1683_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1692_1683_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1684
    process(RPIPE_timer_req_1686_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1686_wire(0 downto 0);
      req_1684 <= tmp_var; -- 
    end process;
    do_while_stmt_1677_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1698_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1677_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1677_branch_req_0,
          ack0 => do_while_stmt_1677_branch_ack_0,
          ack1 => do_while_stmt_1677_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1691_inst
    process(COUNTER_1679) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1679, konst_1690_wire_constant, tmp_var);
      nCOUNTER_1692 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1686_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1686_inst_req_0;
      RPIPE_timer_req_1686_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1686_inst_req_1;
      RPIPE_timer_req_1686_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1686_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1694_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1694_inst_req_0;
      WPIPE_timer_resp_1694_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1694_inst_req_1;
      WPIPE_timer_resp_1694_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1684(0);
      data_in <= COUNTER_1679;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Concat_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    Concat_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    Concat_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module concat
  component concat is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
      Concat_input_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
      Concat_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module concat
  signal concat_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal concat_tag_out   : std_logic_vector(1 downto 0);
  signal concat_start_req : std_logic;
  signal concat_start_ack : std_logic;
  signal concat_fin_req   : std_logic;
  signal concat_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for read from pipe Concat_input_pipe
  signal Concat_input_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal Concat_input_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal Concat_input_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Concat_output_pipe
  signal Concat_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal Concat_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal Concat_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module concat
  concat_instance:concat-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => concat_start_req,
      start_ack => concat_start_ack,
      fin_req => concat_fin_req,
      fin_ack => concat_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      Concat_input_pipe_pipe_read_req => Concat_input_pipe_pipe_read_req(1 downto 0),
      Concat_input_pipe_pipe_read_ack => Concat_input_pipe_pipe_read_ack(1 downto 0),
      Concat_input_pipe_pipe_read_data => Concat_input_pipe_pipe_read_data(15 downto 0),
      Concat_output_pipe_pipe_write_req => Concat_output_pipe_pipe_write_req(0 downto 0),
      Concat_output_pipe_pipe_write_ack => Concat_output_pipe_pipe_write_ack(0 downto 0),
      Concat_output_pipe_pipe_write_data => Concat_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => concat_tag_in,
      tag_out => concat_tag_out-- 
    ); -- 
  -- module will be run forever 
  concat_tag_in <= (others => '0');
  concat_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => concat_start_req, start_ack => concat_start_ack,  fin_req => concat_fin_req,  fin_ack => concat_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  Concat_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_input_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Concat_input_pipe_pipe_read_req,
      read_ack => Concat_input_pipe_pipe_read_ack,
      read_data => Concat_input_pipe_pipe_read_data,
      write_req => Concat_input_pipe_pipe_write_req,
      write_ack => Concat_input_pipe_pipe_write_ack,
      write_data => Concat_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Concat_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Concat_output_pipe_pipe_read_req,
      read_ack => Concat_output_pipe_pipe_read_ack,
      read_data => Concat_output_pipe_pipe_read_data,
      write_req => Concat_output_pipe_pipe_write_req,
      write_ack => Concat_output_pipe_pipe_write_ack,
      write_data => Concat_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
